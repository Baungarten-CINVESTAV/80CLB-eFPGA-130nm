magic
tech sky130A
magscale 1 2
timestamp 1707851634
<< viali >>
rect 6837 9673 6871 9707
rect 2329 9605 2363 9639
rect 3525 9605 3559 9639
rect 4721 9605 4755 9639
rect 9505 9605 9539 9639
rect 1593 9537 1627 9571
rect 1961 9537 1995 9571
rect 2421 9537 2455 9571
rect 2881 9521 2915 9555
rect 3157 9537 3191 9571
rect 4353 9537 4387 9571
rect 5549 9537 5583 9571
rect 6745 9537 6779 9571
rect 7941 9537 7975 9571
rect 8769 9537 8803 9571
rect 9137 9537 9171 9571
rect 9781 9537 9815 9571
rect 10149 9537 10183 9571
rect 2605 9401 2639 9435
rect 5733 9401 5767 9435
rect 8125 9401 8159 9435
rect 10333 9401 10367 9435
rect 1409 9333 1443 9367
rect 2697 9333 2731 9367
rect 8585 9333 8619 9367
rect 9965 9333 9999 9367
rect 1593 9129 1627 9163
rect 2053 9129 2087 9163
rect 4537 9129 4571 9163
rect 9229 9129 9263 9163
rect 10241 9129 10275 9163
rect 2237 8925 2271 8959
rect 4721 8925 4755 8959
rect 6285 8925 6319 8959
rect 9413 8925 9447 8959
rect 1501 8857 1535 8891
rect 9597 8857 9631 8891
rect 9965 8857 9999 8891
rect 10149 8857 10183 8891
rect 6101 8789 6135 8823
rect 8953 8585 8987 8619
rect 9321 8585 9355 8619
rect 10241 8585 10275 8619
rect 9965 8517 9999 8551
rect 1409 8449 1443 8483
rect 5365 8449 5399 8483
rect 8769 8449 8803 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 9873 8449 9907 8483
rect 10149 8449 10183 8483
rect 7665 8381 7699 8415
rect 1593 8313 1627 8347
rect 5181 8313 5215 8347
rect 9045 8313 9079 8347
rect 9597 8313 9631 8347
rect 5457 8041 5491 8075
rect 9505 8041 9539 8075
rect 7849 7973 7883 8007
rect 9965 7973 9999 8007
rect 10333 7973 10367 8007
rect 6745 7905 6779 7939
rect 8125 7905 8159 7939
rect 9597 7905 9631 7939
rect 9781 7905 9815 7939
rect 5365 7837 5399 7871
rect 5641 7837 5675 7871
rect 6561 7837 6595 7871
rect 6653 7837 6687 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 7941 7837 7975 7871
rect 9321 7837 9355 7871
rect 10517 7837 10551 7871
rect 9045 7769 9079 7803
rect 5181 7701 5215 7735
rect 6377 7701 6411 7735
rect 8585 7701 8619 7735
rect 9413 7497 9447 7531
rect 10333 7497 10367 7531
rect 8217 7429 8251 7463
rect 8401 7429 8435 7463
rect 8493 7429 8527 7463
rect 1409 7361 1443 7395
rect 1869 7361 1903 7395
rect 5089 7361 5123 7395
rect 5181 7361 5215 7395
rect 6745 7361 6779 7395
rect 7481 7361 7515 7395
rect 7573 7361 7607 7395
rect 9137 7361 9171 7395
rect 9597 7361 9631 7395
rect 10057 7361 10091 7395
rect 10517 7361 10551 7395
rect 5273 7293 5307 7327
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 6561 7293 6595 7327
rect 7757 7293 7791 7327
rect 9045 7293 9079 7327
rect 1593 7225 1627 7259
rect 4905 7225 4939 7259
rect 7205 7225 7239 7259
rect 9873 7225 9907 7259
rect 1685 7157 1719 7191
rect 5825 7157 5859 7191
rect 7297 7157 7331 7191
rect 9229 7157 9263 7191
rect 7481 6953 7515 6987
rect 6469 6885 6503 6919
rect 8493 6885 8527 6919
rect 5089 6817 5123 6851
rect 6745 6817 6779 6851
rect 7941 6817 7975 6851
rect 1593 6749 1627 6783
rect 2053 6749 2087 6783
rect 2513 6749 2547 6783
rect 2789 6749 2823 6783
rect 3065 6749 3099 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 4997 6749 5031 6783
rect 7389 6749 7423 6783
rect 8953 6749 8987 6783
rect 9209 6749 9243 6783
rect 5356 6681 5390 6715
rect 8042 6681 8076 6715
rect 1685 6613 1719 6647
rect 2145 6613 2179 6647
rect 2329 6613 2363 6647
rect 2605 6613 2639 6647
rect 2881 6613 2915 6647
rect 7297 6613 7331 6647
rect 10333 6613 10367 6647
rect 1593 6409 1627 6443
rect 2697 6409 2731 6443
rect 5457 6409 5491 6443
rect 6009 6409 6043 6443
rect 8769 6409 8803 6443
rect 9045 6409 9079 6443
rect 9321 6409 9355 6443
rect 9689 6409 9723 6443
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 2237 6273 2271 6307
rect 2513 6273 2547 6307
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3157 6297 3191 6331
rect 3617 6273 3651 6307
rect 3801 6273 3835 6307
rect 4068 6273 4102 6307
rect 5641 6273 5675 6307
rect 5741 6271 5775 6305
rect 6193 6273 6227 6307
rect 6561 6273 6595 6307
rect 6828 6273 6862 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 9505 6273 9539 6307
rect 9597 6273 9631 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 8125 6205 8159 6239
rect 1685 6137 1719 6171
rect 2053 6137 2087 6171
rect 2973 6137 3007 6171
rect 3433 6137 3467 6171
rect 8677 6137 8711 6171
rect 2329 6069 2363 6103
rect 3341 6069 3375 6103
rect 5181 6069 5215 6103
rect 5825 6069 5859 6103
rect 7941 6069 7975 6103
rect 9873 6069 9907 6103
rect 10241 6069 10275 6103
rect 2421 5865 2455 5899
rect 6101 5865 6135 5899
rect 7205 5865 7239 5899
rect 7665 5865 7699 5899
rect 9229 5865 9263 5899
rect 2697 5797 2731 5831
rect 2973 5797 3007 5831
rect 3249 5797 3283 5831
rect 5181 5797 5215 5831
rect 5457 5797 5491 5831
rect 6653 5729 6687 5763
rect 7481 5729 7515 5763
rect 8033 5729 8067 5763
rect 9045 5729 9079 5763
rect 9689 5729 9723 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 2329 5661 2363 5695
rect 2605 5661 2639 5695
rect 2881 5661 2915 5695
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 4537 5661 4571 5695
rect 5641 5661 5675 5695
rect 5917 5661 5951 5695
rect 6009 5661 6043 5695
rect 6285 5661 6319 5695
rect 7297 5661 7331 5695
rect 8217 5661 8251 5695
rect 8953 5661 8987 5695
rect 9413 5661 9447 5695
rect 9781 5593 9815 5627
rect 10333 5593 10367 5627
rect 1685 5525 1719 5559
rect 1961 5525 1995 5559
rect 2145 5525 2179 5559
rect 4445 5525 4479 5559
rect 5733 5525 5767 5559
rect 6469 5525 6503 5559
rect 8677 5525 8711 5559
rect 1593 5321 1627 5355
rect 4629 5321 4663 5355
rect 5273 5321 5307 5355
rect 10057 5321 10091 5355
rect 4169 5253 4203 5287
rect 1409 5185 1443 5219
rect 1869 5185 1903 5219
rect 2237 5185 2271 5219
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 4453 5185 4487 5219
rect 4561 5185 4595 5219
rect 4997 5185 5031 5219
rect 5457 5185 5491 5219
rect 6377 5185 6411 5219
rect 8401 5185 8435 5219
rect 8668 5185 8702 5219
rect 9965 5185 9999 5219
rect 2329 5117 2363 5151
rect 3341 5117 3375 5151
rect 3525 5117 3559 5151
rect 3709 5117 3743 5151
rect 5549 5117 5583 5151
rect 5733 5117 5767 5151
rect 1961 5049 1995 5083
rect 4261 5049 4295 5083
rect 5089 5049 5123 5083
rect 6193 5049 6227 5083
rect 2513 4981 2547 5015
rect 2789 4981 2823 5015
rect 7665 4981 7699 5015
rect 9781 4981 9815 5015
rect 4629 4777 4663 4811
rect 9597 4777 9631 4811
rect 3249 4709 3283 4743
rect 5549 4709 5583 4743
rect 6009 4709 6043 4743
rect 6929 4709 6963 4743
rect 8769 4709 8803 4743
rect 2605 4641 2639 4675
rect 4905 4641 4939 4675
rect 6561 4641 6595 4675
rect 7205 4641 7239 4675
rect 9045 4641 9079 4675
rect 9873 4641 9907 4675
rect 10149 4641 10183 4675
rect 1501 4573 1535 4607
rect 2329 4573 2363 4607
rect 2421 4573 2455 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4537 4573 4571 4607
rect 5089 4573 5123 4607
rect 5641 4573 5675 4607
rect 5825 4573 5859 4607
rect 6377 4573 6411 4607
rect 7113 4573 7147 4607
rect 7389 4573 7423 4607
rect 7656 4505 7690 4539
rect 9965 4505 9999 4539
rect 1593 4437 1627 4471
rect 2145 4437 2179 4471
rect 3065 4437 3099 4471
rect 3525 4437 3559 4471
rect 4445 4437 4479 4471
rect 1961 4233 1995 4267
rect 3709 4233 3743 4267
rect 8677 4233 8711 4267
rect 10333 4233 10367 4267
rect 1501 4165 1535 4199
rect 7205 4165 7239 4199
rect 2145 4097 2179 4131
rect 2596 4097 2630 4131
rect 3985 4097 4019 4131
rect 4261 4097 4295 4131
rect 4445 4097 4479 4131
rect 4997 4097 5031 4131
rect 5733 4097 5767 4131
rect 6193 4097 6227 4131
rect 7665 4097 7699 4131
rect 8953 4097 8987 4131
rect 9873 4097 9907 4131
rect 2329 4029 2363 4063
rect 4077 4029 4111 4063
rect 5181 4029 5215 4063
rect 6377 4029 6411 4063
rect 7021 4029 7055 4063
rect 8033 4029 8067 4063
rect 9689 4029 9723 4063
rect 1593 3893 1627 3927
rect 4905 3893 4939 3927
rect 5457 3893 5491 3927
rect 5917 3893 5951 3927
rect 6009 3893 6043 3927
rect 7297 3893 7331 3927
rect 7757 3893 7791 3927
rect 9597 3893 9631 3927
rect 1777 3689 1811 3723
rect 4077 3689 4111 3723
rect 4997 3689 5031 3723
rect 8309 3689 8343 3723
rect 3617 3621 3651 3655
rect 6101 3621 6135 3655
rect 10333 3621 10367 3655
rect 2973 3553 3007 3587
rect 3157 3553 3191 3587
rect 4261 3553 4295 3587
rect 6929 3553 6963 3587
rect 1593 3485 1627 3519
rect 2697 3485 2731 3519
rect 3893 3485 3927 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 4629 3485 4663 3519
rect 5365 3485 5399 3519
rect 6469 3485 6503 3519
rect 7196 3485 7230 3519
rect 8585 3485 8619 3519
rect 2053 3417 2087 3451
rect 2421 3417 2455 3451
rect 5549 3417 5583 3451
rect 5641 3417 5675 3451
rect 9321 3417 9355 3451
rect 9781 3417 9815 3451
rect 9873 3417 9907 3451
rect 2789 3349 2823 3383
rect 5181 3349 5215 3383
rect 6745 3349 6779 3383
rect 8401 3349 8435 3383
rect 2237 3145 2271 3179
rect 9137 3145 9171 3179
rect 10241 3145 10275 3179
rect 1777 3077 1811 3111
rect 2605 3077 2639 3111
rect 4169 3077 4203 3111
rect 4690 3077 4724 3111
rect 7849 3077 7883 3111
rect 9781 3077 9815 3111
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 4445 3009 4479 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6644 3009 6678 3043
rect 10425 3009 10459 3043
rect 2421 2873 2455 2907
rect 7757 2873 7791 2907
rect 5825 2805 5859 2839
rect 6193 2805 6227 2839
rect 9873 2805 9907 2839
rect 8585 2601 8619 2635
rect 2605 2533 2639 2567
rect 2973 2533 3007 2567
rect 7757 2533 7791 2567
rect 8217 2533 8251 2567
rect 9597 2533 9631 2567
rect 2145 2465 2179 2499
rect 2329 2465 2363 2499
rect 3893 2465 3927 2499
rect 6193 2465 6227 2499
rect 7113 2465 7147 2499
rect 7297 2465 7331 2499
rect 7849 2465 7883 2499
rect 8033 2465 8067 2499
rect 9045 2465 9079 2499
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 4261 2397 4295 2431
rect 4997 2397 5031 2431
rect 6653 2397 6687 2431
rect 8769 2397 8803 2431
rect 10333 2397 10367 2431
rect 1685 2329 1719 2363
rect 2053 2329 2087 2363
rect 5549 2329 5583 2363
rect 5641 2329 5675 2363
rect 9137 2329 9171 2363
rect 9873 2329 9907 2363
rect 3341 2261 3375 2295
rect 4353 2261 4387 2295
rect 5089 2261 5123 2295
rect 6929 2261 6963 2295
rect 9965 2261 9999 2295
rect 10517 2261 10551 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6604 9676 6837 9704
rect 6604 9664 6610 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 9582 9704 9588 9716
rect 6825 9667 6883 9673
rect 8772 9676 9588 9704
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 2317 9639 2375 9645
rect 2317 9636 2329 9639
rect 1820 9608 2329 9636
rect 1820 9596 1826 9608
rect 2317 9605 2329 9608
rect 2363 9605 2375 9639
rect 2317 9599 2375 9605
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3513 9639 3571 9645
rect 3513 9636 3525 9639
rect 3016 9608 3525 9636
rect 3016 9596 3022 9608
rect 3513 9605 3525 9608
rect 3559 9605 3571 9639
rect 3513 9599 3571 9605
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4212 9608 4721 9636
rect 4212 9596 4218 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 4709 9599 4767 9605
rect 934 9528 940 9580
rect 992 9568 998 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 992 9540 1593 9568
rect 992 9528 998 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2406 9528 2412 9580
rect 2464 9528 2470 9580
rect 3145 9571 3203 9577
rect 2869 9555 2927 9561
rect 2869 9552 2881 9555
rect 2792 9524 2881 9552
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 2792 9500 2820 9524
rect 2869 9521 2881 9524
rect 2915 9521 2927 9555
rect 3145 9537 3157 9571
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 2869 9515 2927 9521
rect 2740 9472 2820 9500
rect 2740 9460 2746 9472
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3160 9500 3188 9531
rect 4338 9528 4344 9580
rect 4396 9528 4402 9580
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 8772 9577 8800 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 8996 9608 9505 9636
rect 8996 9596 9002 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9784 9608 10548 9636
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 5776 9540 6745 9568
rect 5776 9528 5782 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 3016 9472 3188 9500
rect 7944 9500 7972 9531
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9784 9577 9812 9608
rect 10520 9580 10548 9608
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 7944 9472 9168 9500
rect 3016 9460 3022 9472
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2639 9404 5304 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 1394 9324 1400 9376
rect 1452 9324 1458 9376
rect 2682 9324 2688 9376
rect 2740 9324 2746 9376
rect 5276 9364 5304 9404
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 5721 9435 5779 9441
rect 5721 9432 5733 9435
rect 5408 9404 5733 9432
rect 5408 9392 5414 9404
rect 5721 9401 5733 9404
rect 5767 9401 5779 9435
rect 5721 9395 5779 9401
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 8113 9435 8171 9441
rect 8113 9432 8125 9435
rect 7800 9404 8125 9432
rect 7800 9392 7806 9404
rect 8113 9401 8125 9404
rect 8159 9401 8171 9435
rect 9140 9432 9168 9472
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 10152 9500 10180 9531
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 9272 9472 10180 9500
rect 9272 9460 9278 9472
rect 10042 9432 10048 9444
rect 9140 9404 10048 9432
rect 8113 9395 8171 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 10192 9404 10333 9432
rect 10192 9392 10198 9404
rect 10321 9401 10333 9404
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 7834 9364 7840 9376
rect 5276 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 9030 9364 9036 9376
rect 8619 9336 9036 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9950 9324 9956 9376
rect 10008 9324 10014 9376
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 566 9120 572 9172
rect 624 9160 630 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 624 9132 1593 9160
rect 624 9120 630 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2041 9163 2099 9169
rect 2041 9160 2053 9163
rect 2004 9132 2053 9160
rect 2004 9120 2010 9132
rect 2041 9129 2053 9132
rect 2087 9129 2099 9163
rect 2041 9123 2099 9129
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2740 9120 2774 9160
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4396 9132 4537 9160
rect 4396 9120 4402 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 9214 9120 9220 9172
rect 9272 9120 9278 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9364 9132 10241 9160
rect 9364 9120 9370 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 2746 9024 2774 9120
rect 9950 9052 9956 9104
rect 10008 9052 10014 9104
rect 2746 8996 6316 9024
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2056 8928 2237 8956
rect 1486 8848 1492 8900
rect 1544 8848 1550 8900
rect 2056 8832 2084 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 6288 8965 6316 8996
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4304 8928 4721 8956
rect 4304 8916 4310 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9968 8956 9996 9052
rect 11330 8956 11336 8968
rect 9447 8928 9996 8956
rect 10060 8928 11336 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9582 8848 9588 8900
rect 9640 8848 9646 8900
rect 9953 8891 10011 8897
rect 9953 8857 9965 8891
rect 9999 8888 10011 8891
rect 10060 8888 10088 8928
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 9999 8860 10088 8888
rect 9999 8857 10011 8860
rect 9953 8851 10011 8857
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10192 8860 10237 8888
rect 10192 8848 10198 8860
rect 2038 8780 2044 8832
rect 2096 8780 2102 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 6638 8820 6644 8832
rect 6135 8792 6644 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 9214 8780 9220 8832
rect 9272 8820 9278 8832
rect 10134 8820 10162 8848
rect 9272 8792 10162 8820
rect 9272 8780 9278 8792
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 1394 8576 1400 8628
rect 1452 8576 1458 8628
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 2096 8588 8953 8616
rect 2096 8576 2102 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 9180 8588 9321 8616
rect 9180 8576 9186 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 9640 8588 10241 8616
rect 9640 8576 9646 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 1412 8548 1440 8576
rect 1412 8520 2774 8548
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2746 8480 2774 8520
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 9953 8551 10011 8557
rect 9953 8548 9965 8551
rect 9456 8520 9965 8548
rect 9456 8508 9462 8520
rect 9953 8517 9965 8520
rect 9999 8517 10011 8551
rect 9953 8511 10011 8517
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 2746 8452 5365 8480
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9769 8483 9827 8489
rect 9539 8452 9628 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 7466 8412 7472 8424
rect 5184 8384 7472 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 1762 8344 1768 8356
rect 1627 8316 1768 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 5184 8353 5212 8384
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7650 8372 7656 8424
rect 7708 8372 7714 8424
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8313 5227 8347
rect 5169 8307 5227 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 9600 8353 9628 8452
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9784 8412 9812 8443
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 9950 8412 9956 8424
rect 9784 8384 9956 8412
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 6972 8316 9045 8344
rect 6972 8304 6978 8316
rect 9033 8313 9045 8316
rect 9079 8313 9091 8347
rect 9033 8307 9091 8313
rect 9585 8347 9643 8353
rect 9585 8313 9597 8347
rect 9631 8313 9643 8347
rect 10152 8344 10180 8443
rect 9585 8307 9643 8313
rect 9692 8316 10180 8344
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9692 8276 9720 8316
rect 9272 8248 9720 8276
rect 9272 8236 9278 8248
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5534 8072 5540 8084
rect 5491 8044 5540 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 5684 8044 9505 8072
rect 5684 8032 5690 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 8004 7895 8007
rect 9953 8007 10011 8013
rect 9953 8004 9965 8007
rect 7883 7976 9965 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 6270 7936 6276 7948
rect 5368 7908 6276 7936
rect 5368 7877 5396 7908
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 6779 7908 8125 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5644 7800 5672 7831
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6917 7871 6975 7877
rect 6687 7840 6868 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 5368 7772 5672 7800
rect 5368 7744 5396 7772
rect 6840 7744 6868 7840
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 7055 7840 7205 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 6932 7800 6960 7831
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8220 7868 8248 7976
rect 9953 7973 9965 7976
rect 9999 7973 10011 8007
rect 9953 7967 10011 7973
rect 10321 8007 10379 8013
rect 10321 7973 10333 8007
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9456 7908 9597 7936
rect 9456 7896 9462 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 10336 7936 10364 7967
rect 9815 7908 10364 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 7975 7840 8248 7868
rect 8956 7840 9321 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8956 7800 8984 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10008 7840 10517 7868
rect 10008 7828 10014 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 6932 7772 7880 7800
rect 7852 7744 7880 7772
rect 8128 7772 8984 7800
rect 9033 7803 9091 7809
rect 8128 7744 8156 7772
rect 9033 7769 9045 7803
rect 9079 7800 9091 7803
rect 9858 7800 9864 7812
rect 9079 7772 9864 7800
rect 9079 7769 9091 7772
rect 9033 7763 9091 7769
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 6362 7692 6368 7744
rect 6420 7692 6426 7744
rect 6822 7692 6828 7744
rect 6880 7692 6886 7744
rect 7834 7692 7840 7744
rect 7892 7692 7898 7744
rect 8110 7692 8116 7744
rect 8168 7692 8174 7744
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 8662 7732 8668 7744
rect 8619 7704 8668 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 6362 7488 6368 7540
rect 6420 7488 6426 7540
rect 8662 7528 8668 7540
rect 8404 7500 8668 7528
rect 5184 7460 5212 7488
rect 5092 7432 5212 7460
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1854 7352 1860 7404
rect 1912 7352 1918 7404
rect 5092 7401 5120 7432
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5350 7392 5356 7404
rect 5215 7364 5356 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 5184 7324 5212 7355
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6380 7392 6408 7488
rect 8404 7469 8432 7500
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9950 7528 9956 7540
rect 9447 7500 9956 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10321 7531 10379 7537
rect 10321 7497 10333 7531
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7460 8263 7463
rect 8389 7463 8447 7469
rect 8389 7460 8401 7463
rect 8251 7432 8401 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 8389 7429 8401 7432
rect 8435 7429 8447 7463
rect 8389 7423 8447 7429
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7460 8539 7463
rect 9306 7460 9312 7472
rect 8527 7432 9312 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6380 7364 6745 7392
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 6880 7364 7481 7392
rect 6880 7352 6886 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7650 7392 7656 7404
rect 7607 7364 7656 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9456 7364 9597 7392
rect 9456 7352 9462 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10336 7392 10364 7491
rect 10091 7364 10364 7392
rect 10505 7395 10563 7401
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10870 7392 10876 7404
rect 10551 7364 10876 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 1544 7296 5212 7324
rect 5261 7327 5319 7333
rect 1544 7284 1550 7296
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5307 7296 5457 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 5629 7287 5687 7293
rect 5828 7296 6561 7324
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2498 7256 2504 7268
rect 1627 7228 2504 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5644 7256 5672 7287
rect 4939 7228 5672 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5828 7200 5856 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 7742 7284 7748 7336
rect 7800 7284 7806 7336
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9232 7324 9260 7352
rect 9079 7296 9260 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 7193 7259 7251 7265
rect 7193 7225 7205 7259
rect 7239 7256 7251 7259
rect 7650 7256 7656 7268
rect 7239 7228 7656 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 9861 7259 9919 7265
rect 7892 7228 9352 7256
rect 7892 7216 7898 7228
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 2866 7188 2872 7200
rect 1719 7160 2872 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 5810 7148 5816 7200
rect 5868 7148 5874 7200
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 8662 7188 8668 7200
rect 7331 7160 8668 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8904 7160 9229 7188
rect 8904 7148 8910 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9324 7188 9352 7228
rect 9861 7225 9873 7259
rect 9907 7256 9919 7259
rect 10042 7256 10048 7268
rect 9907 7228 10048 7256
rect 9907 7225 9919 7228
rect 9861 7219 9919 7225
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10410 7188 10416 7200
rect 9324 7160 10416 7188
rect 9217 7151 9275 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2372 6956 7328 6984
rect 2372 6944 2378 6956
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 2556 6888 3372 6916
rect 2556 6876 2562 6888
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 1596 6712 1624 6743
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1912 6752 2053 6780
rect 1912 6740 1918 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 2516 6712 2544 6743
rect 2774 6740 2780 6792
rect 2832 6740 2838 6792
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3344 6780 3372 6888
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 6512 6888 6776 6916
rect 6512 6876 6518 6888
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 6748 6857 6776 6888
rect 7300 6860 7328 6956
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7432 6956 7481 6984
rect 7432 6944 7438 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 9214 6984 9220 6996
rect 7469 6947 7527 6953
rect 8496 6956 9220 6984
rect 7650 6876 7656 6928
rect 7708 6876 7714 6928
rect 8496 6925 8524 6956
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 8481 6919 8539 6925
rect 8481 6885 8493 6919
rect 8527 6885 8539 6919
rect 8481 6879 8539 6885
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 3936 6820 5089 6848
rect 3936 6808 3942 6820
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 6822 6848 6828 6860
rect 6779 6820 6828 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7282 6808 7288 6860
rect 7340 6808 7346 6860
rect 7668 6848 7696 6876
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7668 6820 7941 6848
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3344 6752 4077 6780
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4203 6752 4353 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5810 6780 5816 6792
rect 5031 6752 5816 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 3234 6712 3240 6724
rect 1596 6684 3240 6712
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 1670 6604 1676 6656
rect 1728 6604 1734 6656
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 2004 6616 2145 6644
rect 2004 6604 2010 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2498 6644 2504 6656
rect 2363 6616 2504 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2590 6604 2596 6656
rect 2648 6604 2654 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3694 6644 3700 6656
rect 2915 6616 3700 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4540 6644 4568 6743
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 6328 6752 7389 6780
rect 6328 6740 6334 6752
rect 7377 6749 7389 6752
rect 7423 6780 7435 6783
rect 7423 6752 7604 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 5344 6715 5402 6721
rect 5344 6681 5356 6715
rect 5390 6712 5402 6715
rect 6362 6712 6368 6724
rect 5390 6684 6368 6712
rect 5390 6681 5402 6684
rect 5344 6675 5402 6681
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 7576 6656 7604 6752
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9197 6783 9255 6789
rect 9197 6780 9209 6783
rect 9088 6752 9209 6780
rect 9088 6740 9094 6752
rect 9197 6749 9209 6752
rect 9243 6749 9255 6783
rect 9197 6743 9255 6749
rect 8030 6715 8088 6721
rect 8030 6681 8042 6715
rect 8076 6712 8088 6715
rect 8076 6684 8156 6712
rect 8076 6681 8088 6684
rect 8030 6675 8088 6681
rect 6178 6644 6184 6656
rect 4540 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 8128 6644 8156 6684
rect 9398 6672 9404 6724
rect 9456 6712 9462 6724
rect 9456 6684 10364 6712
rect 9456 6672 9462 6684
rect 9674 6644 9680 6656
rect 8128 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10336 6653 10364 6684
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1627 6412 1900 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1762 6332 1768 6384
rect 1820 6332 1826 6384
rect 1872 6372 1900 6412
rect 2314 6400 2320 6452
rect 2372 6400 2378 6452
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 3050 6440 3056 6452
rect 2731 6412 3056 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 5166 6440 5172 6452
rect 3252 6412 5172 6440
rect 2332 6372 2360 6400
rect 1872 6344 2360 6372
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1780 6236 1808 6332
rect 1872 6313 1900 6344
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2424 6304 2452 6400
rect 2700 6344 3096 6372
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 2424 6276 2513 6304
rect 2225 6267 2283 6273
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2240 6236 2268 6267
rect 1780 6208 2268 6236
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 2608 6236 2636 6267
rect 2464 6208 2636 6236
rect 2464 6196 2470 6208
rect 1670 6128 1676 6180
rect 1728 6128 1734 6180
rect 2041 6171 2099 6177
rect 2041 6137 2053 6171
rect 2087 6168 2099 6171
rect 2700 6168 2728 6344
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 2087 6140 2728 6168
rect 2087 6137 2099 6140
rect 2041 6131 2099 6137
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 1636 6072 2329 6100
rect 1636 6060 1642 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2884 6100 2912 6267
rect 3068 6236 3096 6344
rect 3160 6337 3188 6400
rect 3145 6331 3203 6337
rect 3145 6297 3157 6331
rect 3191 6297 3203 6331
rect 3145 6291 3203 6297
rect 3252 6236 3280 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6440 5503 6443
rect 5718 6440 5724 6452
rect 5491 6412 5724 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6546 6440 6552 6452
rect 6043 6412 6552 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 7800 6412 8769 6440
rect 7800 6400 7806 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 8938 6400 8944 6452
rect 8996 6400 9002 6452
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 4982 6332 4988 6384
rect 5040 6372 5046 6384
rect 5534 6372 5540 6384
rect 5040 6344 5540 6372
rect 5040 6332 5046 6344
rect 5534 6332 5540 6344
rect 5592 6372 5598 6384
rect 5592 6344 5672 6372
rect 5592 6332 5598 6344
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 3878 6304 3884 6316
rect 3835 6276 3884 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 5644 6313 5672 6344
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 6270 6372 6276 6384
rect 6144 6344 6276 6372
rect 6144 6332 6150 6344
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 6454 6332 6460 6384
rect 6512 6332 6518 6384
rect 8956 6372 8984 6400
rect 6564 6344 8984 6372
rect 4056 6307 4114 6313
rect 4056 6273 4068 6307
rect 4102 6304 4114 6307
rect 5629 6307 5687 6313
rect 4102 6276 5488 6304
rect 4102 6273 4114 6276
rect 4056 6267 4114 6273
rect 3068 6208 3280 6236
rect 5460 6236 5488 6276
rect 5629 6273 5641 6307
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5729 6305 5787 6311
rect 5729 6271 5741 6305
rect 5775 6302 5787 6305
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 5828 6302 6193 6304
rect 5775 6276 6193 6302
rect 5775 6274 5856 6276
rect 5775 6271 5787 6274
rect 5729 6265 5787 6271
rect 6181 6273 6193 6276
rect 6227 6304 6239 6307
rect 6472 6304 6500 6332
rect 6564 6313 6592 6344
rect 6227 6276 6500 6304
rect 6549 6307 6607 6313
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6816 6307 6874 6313
rect 6816 6273 6828 6307
rect 6862 6304 6874 6307
rect 7282 6304 7288 6316
rect 6862 6276 7288 6304
rect 6862 6273 6874 6276
rect 6816 6267 6874 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8720 6276 8953 6304
rect 8720 6264 8726 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 6270 6236 6276 6248
rect 5460 6208 6276 6236
rect 6270 6196 6276 6208
rect 6328 6196 6334 6248
rect 6362 6196 6368 6248
rect 6420 6196 6426 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7616 6208 8125 6236
rect 7616 6196 7622 6208
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 9048 6236 9076 6403
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 9232 6344 9628 6372
rect 9232 6316 9260 6344
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9600 6313 9628 6344
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9508 6236 9536 6267
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10318 6304 10324 6316
rect 10183 6276 10324 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 8159 6208 8800 6236
rect 9048 6208 9536 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 2961 6171 3019 6177
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 3142 6168 3148 6180
rect 3007 6140 3148 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3421 6171 3479 6177
rect 3421 6137 3433 6171
rect 3467 6168 3479 6171
rect 3510 6168 3516 6180
rect 3467 6140 3516 6168
rect 3467 6137 3479 6140
rect 3421 6131 3479 6137
rect 3510 6128 3516 6140
rect 3568 6128 3574 6180
rect 3234 6100 3240 6112
rect 2884 6072 3240 6100
rect 2317 6063 2375 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3329 6103 3387 6109
rect 3329 6069 3341 6103
rect 3375 6100 3387 6103
rect 3694 6100 3700 6112
rect 3375 6072 3700 6100
rect 3375 6069 3387 6072
rect 3329 6063 3387 6069
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4488 6072 5181 6100
rect 4488 6060 4494 6072
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 5169 6063 5227 6069
rect 5810 6060 5816 6112
rect 5868 6060 5874 6112
rect 6380 6100 6408 6196
rect 8665 6171 8723 6177
rect 8665 6168 8677 6171
rect 7484 6140 8677 6168
rect 7484 6100 7512 6140
rect 8665 6137 8677 6140
rect 8711 6137 8723 6171
rect 8772 6168 8800 6208
rect 9398 6168 9404 6180
rect 8772 6140 9404 6168
rect 8665 6131 8723 6137
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 6380 6072 7512 6100
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7892 6072 7941 6100
rect 7892 6060 7898 6072
rect 7929 6069 7941 6072
rect 7975 6100 7987 6103
rect 9214 6100 9220 6112
rect 7975 6072 9220 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9858 6060 9864 6112
rect 9916 6060 9922 6112
rect 10226 6060 10232 6112
rect 10284 6060 10290 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2774 5896 2780 5908
rect 2455 5868 2780 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 4430 5896 4436 5908
rect 2884 5868 4436 5896
rect 1872 5760 1900 5856
rect 2685 5831 2743 5837
rect 2685 5797 2697 5831
rect 2731 5828 2743 5831
rect 2884 5828 2912 5868
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 6089 5899 6147 5905
rect 5132 5868 5856 5896
rect 5132 5856 5138 5868
rect 2731 5800 2912 5828
rect 2961 5831 3019 5837
rect 2731 5797 2743 5800
rect 2685 5791 2743 5797
rect 2961 5797 2973 5831
rect 3007 5797 3019 5831
rect 2961 5791 3019 5797
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 3283 5800 3924 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 2976 5760 3004 5791
rect 1872 5732 2728 5760
rect 2976 5732 3464 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2038 5692 2044 5704
rect 1903 5664 2044 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1596 5624 1624 5655
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2700 5692 2728 5732
rect 2774 5692 2780 5704
rect 2639 5664 2780 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3326 5692 3332 5704
rect 3191 5664 3332 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3436 5701 3464 5732
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 3896 5692 3924 5800
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 5169 5831 5227 5837
rect 5169 5828 5181 5831
rect 4120 5800 5181 5828
rect 4120 5788 4126 5800
rect 5169 5797 5181 5800
rect 5215 5797 5227 5831
rect 5169 5791 5227 5797
rect 5445 5831 5503 5837
rect 5445 5797 5457 5831
rect 5491 5828 5503 5831
rect 5718 5828 5724 5840
rect 5491 5800 5724 5828
rect 5491 5797 5503 5800
rect 5445 5791 5503 5797
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 5828 5760 5856 5868
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6178 5896 6184 5908
rect 6135 5868 6184 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6328 5868 7205 5896
rect 6328 5856 6334 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 8846 5896 8852 5908
rect 7944 5868 8852 5896
rect 7834 5828 7840 5840
rect 6656 5800 7840 5828
rect 6086 5760 6092 5772
rect 5828 5732 6092 5760
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3896 5664 3985 5692
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 4338 5692 4344 5704
rect 3973 5655 4031 5661
rect 4071 5664 4344 5692
rect 3344 5624 3372 5652
rect 4071 5624 4099 5664
rect 4338 5652 4344 5664
rect 4396 5692 4402 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4396 5664 4537 5692
rect 4396 5652 4402 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6012 5701 6040 5732
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6656 5769 6684 5800
rect 7834 5788 7840 5800
rect 7892 5788 7898 5840
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 7469 5763 7527 5769
rect 7469 5760 7481 5763
rect 6788 5732 7481 5760
rect 6788 5720 6794 5732
rect 7469 5729 7481 5732
rect 7515 5729 7527 5763
rect 7469 5723 7527 5729
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 5592 5664 5641 5692
rect 5592 5652 5598 5664
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5951 5664 6009 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5692 6331 5695
rect 6822 5692 6828 5704
rect 6319 5664 6828 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6972 5664 7297 5692
rect 6972 5652 6978 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7944 5692 7972 5868
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 10042 5896 10048 5908
rect 9263 5868 10048 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 9950 5828 9956 5840
rect 9692 5800 9956 5828
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8067 5732 9045 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9692 5769 9720 5800
rect 9950 5788 9956 5800
rect 10008 5788 10014 5840
rect 9677 5763 9735 5769
rect 9180 5732 9444 5760
rect 9180 5720 9186 5732
rect 9416 5701 9444 5732
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7944 5664 8217 5692
rect 7285 5655 7343 5661
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8205 5655 8263 5661
rect 8312 5664 8953 5692
rect 6178 5624 6184 5636
rect 1596 5596 2820 5624
rect 3344 5596 4099 5624
rect 4172 5596 6184 5624
rect 1670 5516 1676 5568
rect 1728 5516 1734 5568
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2038 5556 2044 5568
rect 1995 5528 2044 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 2682 5556 2688 5568
rect 2179 5528 2688 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 2792 5556 2820 5596
rect 4172 5568 4200 5596
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 8110 5624 8116 5636
rect 6472 5596 8116 5624
rect 2866 5556 2872 5568
rect 2792 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5556 2930 5568
rect 3694 5556 3700 5568
rect 2924 5528 3700 5556
rect 2924 5516 2930 5528
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4706 5556 4712 5568
rect 4479 5528 4712 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6472 5565 6500 5596
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5684 5528 5733 5556
rect 5684 5516 5690 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5525 6515 5559
rect 6457 5519 6515 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 8312 5556 8340 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 8444 5596 9781 5624
rect 8444 5584 8450 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 9950 5584 9956 5636
rect 10008 5624 10014 5636
rect 10321 5627 10379 5633
rect 10321 5624 10333 5627
rect 10008 5596 10333 5624
rect 10008 5584 10014 5596
rect 10321 5593 10333 5596
rect 10367 5593 10379 5627
rect 10321 5587 10379 5593
rect 7432 5528 8340 5556
rect 8665 5559 8723 5565
rect 7432 5516 7438 5528
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 9398 5556 9404 5568
rect 8711 5528 9404 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1596 5284 1624 5315
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1820 5324 3280 5352
rect 1820 5312 1826 5324
rect 1596 5256 2268 5284
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1854 5176 1860 5228
rect 1912 5176 1918 5228
rect 2240 5225 2268 5256
rect 2866 5244 2872 5296
rect 2924 5244 2930 5296
rect 3142 5244 3148 5296
rect 3200 5244 3206 5296
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2271 5188 2697 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2884 5216 2912 5244
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2884 5188 2973 5216
rect 2685 5179 2743 5185
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 3050 5148 3056 5160
rect 2363 5120 3056 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3160 5148 3188 5244
rect 3252 5225 3280 5324
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 3844 5324 4629 5352
rect 3844 5312 3850 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 4706 5312 4712 5364
rect 4764 5312 4770 5364
rect 4890 5312 4896 5364
rect 4948 5312 4954 5364
rect 5074 5352 5080 5364
rect 5000 5324 5080 5352
rect 4157 5287 4215 5293
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4724 5284 4752 5312
rect 4203 5256 4752 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4264 5228 4292 5256
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 4246 5176 4252 5228
rect 4304 5176 4310 5228
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4441 5219 4499 5225
rect 4441 5216 4453 5219
rect 4396 5188 4453 5216
rect 4396 5176 4402 5188
rect 4441 5185 4453 5188
rect 4487 5185 4499 5219
rect 4441 5179 4499 5185
rect 4549 5219 4607 5225
rect 4549 5185 4561 5219
rect 4595 5216 4607 5219
rect 4908 5216 4936 5312
rect 5000 5225 5028 5324
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 6086 5352 6092 5364
rect 5307 5324 6092 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 8812 5324 10057 5352
rect 8812 5312 8818 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 8404 5256 8984 5284
rect 8404 5228 8432 5256
rect 8956 5228 8984 5256
rect 4595 5188 4936 5216
rect 4985 5219 5043 5225
rect 4595 5185 4607 5188
rect 4549 5179 4607 5185
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5626 5216 5632 5228
rect 5491 5188 5632 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 6730 5216 6736 5228
rect 6411 5188 6736 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8662 5225 8668 5228
rect 8656 5179 8668 5225
rect 8662 5176 8668 5179
rect 8720 5176 8726 5228
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9416 5188 9965 5216
rect 3329 5151 3387 5157
rect 3160 5120 3280 5148
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5080 2007 5083
rect 3142 5080 3148 5092
rect 1995 5052 3148 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 1820 4984 2513 5012
rect 1820 4972 1826 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 2774 4972 2780 5024
rect 2832 4972 2838 5024
rect 3252 5012 3280 5120
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3375 5120 3525 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 3694 5108 3700 5160
rect 3752 5108 3758 5160
rect 5368 5148 5396 5176
rect 4908 5120 5396 5148
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 4908 5080 4936 5120
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 4295 5052 4936 5080
rect 5077 5083 5135 5089
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 5077 5049 5089 5083
rect 5123 5080 5135 5083
rect 5736 5080 5764 5111
rect 5123 5052 5764 5080
rect 6181 5083 6239 5089
rect 5123 5049 5135 5052
rect 5077 5043 5135 5049
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6914 5080 6920 5092
rect 6227 5052 6920 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7576 5052 8432 5080
rect 7576 5012 7604 5052
rect 3252 4984 7604 5012
rect 7650 4972 7656 5024
rect 7708 4972 7714 5024
rect 8404 5012 8432 5052
rect 9416 5012 9444 5188
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 8404 4984 9444 5012
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 10134 5012 10140 5024
rect 9815 4984 10140 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 2774 4808 2780 4820
rect 2746 4768 2780 4808
rect 2832 4768 2838 4820
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 3752 4780 4629 4808
rect 3752 4768 3758 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 5460 4780 8616 4808
rect 2746 4740 2774 4768
rect 1504 4712 2774 4740
rect 1504 4613 1532 4712
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2593 4675 2651 4681
rect 2593 4672 2605 4675
rect 2004 4644 2605 4672
rect 2004 4632 2010 4644
rect 2593 4641 2605 4644
rect 2639 4641 2651 4675
rect 2593 4635 2651 4641
rect 2866 4632 2872 4684
rect 2924 4632 2930 4684
rect 3160 4672 3188 4768
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 5460 4740 5488 4780
rect 3283 4712 5488 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 5997 4743 6055 4749
rect 5997 4740 6009 4743
rect 5592 4712 6009 4740
rect 5592 4700 5598 4712
rect 5997 4709 6009 4712
rect 6043 4709 6055 4743
rect 5997 4703 6055 4709
rect 6086 4700 6092 4752
rect 6144 4700 6150 4752
rect 6914 4700 6920 4752
rect 6972 4700 6978 4752
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 3160 4644 4905 4672
rect 4893 4641 4905 4644
rect 4939 4672 4951 4675
rect 6104 4672 6132 4700
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 4939 4644 5212 4672
rect 6104 4644 6561 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 2038 4564 2044 4616
rect 2096 4564 2102 4616
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 2280 4576 2329 4604
rect 2280 4564 2286 4576
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 2056 4536 2084 4564
rect 2424 4536 2452 4567
rect 2056 4508 2452 4536
rect 2884 4536 2912 4632
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 3108 4576 3157 4604
rect 3108 4564 3114 4576
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3145 4567 3203 4573
rect 3344 4576 3433 4604
rect 3344 4536 3372 4576
rect 3421 4573 3433 4576
rect 3467 4604 3479 4607
rect 3786 4604 3792 4616
rect 3467 4576 3792 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4396 4576 4537 4604
rect 4396 4564 4402 4576
rect 4525 4573 4537 4576
rect 4571 4604 4583 4607
rect 4614 4604 4620 4616
rect 4571 4576 4620 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5074 4564 5080 4616
rect 5132 4564 5138 4616
rect 5184 4604 5212 4644
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 6549 4635 6607 4641
rect 6656 4644 7205 4672
rect 5442 4604 5448 4616
rect 5184 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5644 4536 5672 4567
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5776 4576 5825 4604
rect 5776 4564 5782 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6656 4604 6684 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 8386 4632 8392 4684
rect 8444 4632 8450 4684
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6411 4576 6684 4604
rect 6840 4576 7113 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6380 4536 6408 4567
rect 6840 4548 6868 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 8404 4604 8432 4632
rect 7423 4576 8432 4604
rect 8588 4604 8616 4780
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 8720 4780 9597 4808
rect 8720 4768 8726 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4709 8815 4743
rect 8757 4703 8815 4709
rect 8772 4672 8800 4703
rect 9398 4700 9404 4752
rect 9456 4740 9462 4752
rect 9456 4712 9904 4740
rect 9456 4700 9462 4712
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8772 4644 9045 4672
rect 9033 4641 9045 4644
rect 9079 4672 9091 4675
rect 9122 4672 9128 4684
rect 9079 4644 9128 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9876 4681 9904 4712
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 10008 4712 10180 4740
rect 10008 4700 10014 4712
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 10042 4672 10048 4684
rect 9907 4644 10048 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10152 4681 10180 4712
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 8588 4576 8800 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 2884 4508 3372 4536
rect 3436 4508 4660 4536
rect 5644 4508 6408 4536
rect 1302 4428 1308 4480
rect 1360 4468 1366 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 1360 4440 1593 4468
rect 1360 4428 1366 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 2130 4428 2136 4480
rect 2188 4428 2194 4480
rect 3050 4428 3056 4480
rect 3108 4428 3114 4480
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3436 4468 3464 4508
rect 3200 4440 3464 4468
rect 3513 4471 3571 4477
rect 3200 4428 3206 4440
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 4338 4468 4344 4480
rect 3559 4440 4344 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 4522 4468 4528 4480
rect 4479 4440 4528 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4632 4468 4660 4508
rect 6822 4496 6828 4548
rect 6880 4496 6886 4548
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7392 4536 7420 4567
rect 6972 4508 7420 4536
rect 7644 4539 7702 4545
rect 6972 4496 6978 4508
rect 7644 4505 7656 4539
rect 7690 4536 7702 4539
rect 8662 4536 8668 4548
rect 7690 4508 8668 4536
rect 7690 4505 7702 4508
rect 7644 4499 7702 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 8772 4536 8800 4576
rect 9953 4539 10011 4545
rect 8772 4508 9812 4536
rect 7374 4468 7380 4480
rect 4632 4440 7380 4468
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 9784 4468 9812 4508
rect 9953 4505 9965 4539
rect 9999 4505 10011 4539
rect 9953 4499 10011 4505
rect 9968 4468 9996 4499
rect 9784 4440 9996 4468
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1946 4224 1952 4276
rect 2004 4224 2010 4276
rect 2130 4224 2136 4276
rect 2188 4224 2194 4276
rect 3697 4267 3755 4273
rect 3697 4233 3709 4267
rect 3743 4264 3755 4267
rect 3786 4264 3792 4276
rect 3743 4236 3792 4264
rect 3743 4233 3755 4236
rect 3697 4227 3755 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4062 4224 4068 4276
rect 4120 4224 4126 4276
rect 4614 4264 4620 4276
rect 4172 4236 4620 4264
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4196 1547 4199
rect 2148 4196 2176 4224
rect 4080 4196 4108 4224
rect 1535 4168 2176 4196
rect 3896 4168 4108 4196
rect 1535 4165 1547 4168
rect 1489 4159 1547 4165
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2406 4128 2412 4140
rect 2179 4100 2412 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2584 4131 2642 4137
rect 2584 4097 2596 4131
rect 2630 4128 2642 4131
rect 3896 4128 3924 4168
rect 2630 4100 3924 4128
rect 3973 4131 4031 4137
rect 2630 4097 2642 4100
rect 2584 4091 2642 4097
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4172 4128 4200 4236
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 5074 4264 5080 4276
rect 4724 4236 5080 4264
rect 4724 4196 4752 4236
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 5644 4236 8616 4264
rect 5644 4196 5672 4236
rect 6822 4196 6828 4208
rect 4356 4168 4752 4196
rect 4908 4168 5672 4196
rect 5736 4168 6828 4196
rect 4019 4100 4200 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4029 2375 4063
rect 2317 4023 2375 4029
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4060 4123 4063
rect 4356 4060 4384 4168
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 4479 4100 4721 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4111 4032 4384 4060
rect 4693 4060 4721 4100
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 4908 4128 4936 4168
rect 4856 4100 4936 4128
rect 4985 4131 5043 4137
rect 4856 4088 4862 4100
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5534 4128 5540 4140
rect 5031 4100 5540 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5736 4137 5764 4168
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 7193 4199 7251 4205
rect 7193 4165 7205 4199
rect 7239 4196 7251 4199
rect 7466 4196 7472 4208
rect 7239 4168 7472 4196
rect 7239 4165 7251 4168
rect 7193 4159 7251 4165
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 8588 4196 8616 4236
rect 8662 4224 8668 4276
rect 8720 4224 8726 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 10100 4236 10333 4264
rect 10100 4224 10106 4236
rect 10321 4233 10333 4236
rect 10367 4233 10379 4267
rect 10321 4227 10379 4233
rect 9950 4196 9956 4208
rect 8588 4168 9956 4196
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 6227 4100 7665 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 7653 4097 7665 4100
rect 7699 4128 7711 4131
rect 8110 4128 8116 4140
rect 7699 4100 8116 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 8110 4088 8116 4100
rect 8168 4128 8174 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8168 4100 8953 4128
rect 8168 4088 8174 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 4890 4060 4896 4072
rect 4693 4032 4896 4060
rect 4111 4029 4123 4032
rect 4065 4023 4123 4029
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 1946 3992 1952 4004
rect 1728 3964 1952 3992
rect 1728 3952 1734 3964
rect 1946 3952 1952 3964
rect 2004 3952 2010 4004
rect 382 3884 388 3936
rect 440 3924 446 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 440 3896 1593 3924
rect 440 3884 446 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 2332 3924 2360 4023
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 3620 3964 3924 3992
rect 3620 3924 3648 3964
rect 3896 3936 3924 3964
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 5184 3992 5212 4023
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5316 4032 6377 4060
rect 5316 4020 5322 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7466 4060 7472 4072
rect 7055 4032 7472 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 9950 4060 9956 4072
rect 9723 4032 9956 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 4028 3964 5212 3992
rect 4028 3952 4034 3964
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 6328 3964 7328 3992
rect 6328 3952 6334 3964
rect 2332 3896 3648 3924
rect 1581 3887 1639 3893
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4798 3924 4804 3936
rect 4396 3896 4804 3924
rect 4396 3884 4402 3896
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 4982 3924 4988 3936
rect 4939 3896 4988 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5684 3896 5917 3924
rect 5684 3884 5690 3896
rect 5905 3893 5917 3896
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6362 3924 6368 3936
rect 6043 3896 6368 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 7300 3933 7328 3964
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3893 7343 3927
rect 7285 3887 7343 3893
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 7984 3896 9597 3924
rect 7984 3884 7990 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9585 3887 9643 3893
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 1765 3723 1823 3729
rect 1765 3689 1777 3723
rect 1811 3720 1823 3723
rect 2038 3720 2044 3732
rect 1811 3692 2044 3720
rect 1811 3689 1823 3692
rect 1765 3683 1823 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 3050 3720 3056 3732
rect 2700 3692 3056 3720
rect 2590 3544 2596 3596
rect 2648 3584 2654 3596
rect 2700 3584 2728 3692
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 4065 3723 4123 3729
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 4154 3720 4160 3732
rect 4111 3692 4160 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4614 3720 4620 3732
rect 4488 3692 4620 3720
rect 4488 3680 4494 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5534 3720 5540 3732
rect 5040 3692 5540 3720
rect 5040 3680 5046 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6914 3680 6920 3732
rect 6972 3680 6978 3732
rect 7926 3680 7932 3732
rect 7984 3680 7990 3732
rect 8018 3680 8024 3732
rect 8076 3720 8082 3732
rect 8297 3723 8355 3729
rect 8297 3720 8309 3723
rect 8076 3692 8309 3720
rect 8076 3680 8082 3692
rect 8297 3689 8309 3692
rect 8343 3689 8355 3723
rect 8297 3683 8355 3689
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 3605 3655 3663 3661
rect 2832 3624 3188 3652
rect 2832 3612 2838 3624
rect 3160 3593 3188 3624
rect 3605 3621 3617 3655
rect 3651 3652 3663 3655
rect 5442 3652 5448 3664
rect 3651 3624 5448 3652
rect 3651 3621 3663 3624
rect 3605 3615 3663 3621
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 6089 3655 6147 3661
rect 6089 3621 6101 3655
rect 6135 3652 6147 3655
rect 6178 3652 6184 3664
rect 6135 3624 6184 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 6932 3593 6960 3680
rect 2961 3587 3019 3593
rect 2961 3584 2973 3587
rect 2648 3556 2973 3584
rect 2648 3544 2654 3556
rect 2961 3553 2973 3556
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 6917 3587 6975 3593
rect 4295 3556 6500 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1596 3392 1624 3479
rect 2682 3476 2688 3528
rect 2740 3476 2746 3528
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4338 3516 4344 3528
rect 4203 3488 4344 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 2041 3451 2099 3457
rect 2041 3417 2053 3451
rect 2087 3448 2099 3451
rect 2406 3448 2412 3460
rect 2087 3420 2412 3448
rect 2087 3417 2099 3420
rect 2041 3411 2099 3417
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 3510 3408 3516 3460
rect 3568 3408 3574 3460
rect 3896 3448 3924 3479
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4614 3476 4620 3528
rect 4672 3476 4678 3528
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 6472 3525 6500 3556
rect 6917 3553 6929 3587
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 7184 3519 7242 3525
rect 7184 3485 7196 3519
rect 7230 3516 7242 3519
rect 7944 3516 7972 3680
rect 8312 3584 8340 3683
rect 10318 3612 10324 3664
rect 10376 3612 10382 3664
rect 8312 3556 8616 3584
rect 8588 3525 8616 3556
rect 7230 3488 7972 3516
rect 8573 3519 8631 3525
rect 7230 3485 7242 3488
rect 7184 3479 7242 3485
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 5092 3448 5120 3476
rect 3896 3420 5120 3448
rect 5537 3451 5595 3457
rect 5537 3417 5549 3451
rect 5583 3417 5595 3451
rect 5537 3411 5595 3417
rect 5629 3451 5687 3457
rect 5629 3417 5641 3451
rect 5675 3448 5687 3451
rect 5718 3448 5724 3460
rect 5675 3420 5724 3448
rect 5675 3417 5687 3420
rect 5629 3411 5687 3417
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 3528 3380 3556 3408
rect 5169 3383 5227 3389
rect 5169 3380 5181 3383
rect 3528 3352 5181 3380
rect 5169 3349 5181 3352
rect 5215 3349 5227 3383
rect 5169 3343 5227 3349
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5552 3380 5580 3411
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 7668 3420 9321 3448
rect 5500 3352 5580 3380
rect 6733 3383 6791 3389
rect 5500 3340 5506 3352
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7190 3380 7196 3392
rect 6779 3352 7196 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 7668 3380 7696 3420
rect 9309 3417 9321 3420
rect 9355 3448 9367 3451
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 9355 3420 9781 3448
rect 9355 3417 9367 3420
rect 9309 3411 9367 3417
rect 9769 3417 9781 3420
rect 9815 3417 9827 3451
rect 9769 3411 9827 3417
rect 9858 3408 9864 3460
rect 9916 3408 9922 3460
rect 7340 3352 7696 3380
rect 8389 3383 8447 3389
rect 7340 3340 7346 3352
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 9030 3380 9036 3392
rect 8435 3352 9036 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 1452 3148 2237 3176
rect 1452 3136 1458 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 2498 3136 2504 3188
rect 2556 3136 2562 3188
rect 7650 3176 7656 3188
rect 2746 3148 7656 3176
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 2516 3108 2544 3136
rect 1811 3080 2544 3108
rect 2593 3111 2651 3117
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 2056 3049 2084 3080
rect 2593 3077 2605 3111
rect 2639 3108 2651 3111
rect 2746 3108 2774 3148
rect 7650 3136 7656 3148
rect 7708 3176 7714 3188
rect 7708 3148 7880 3176
rect 7708 3136 7714 3148
rect 2639 3080 2774 3108
rect 2639 3077 2651 3080
rect 2593 3071 2651 3077
rect 3878 3068 3884 3120
rect 3936 3108 3942 3120
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 3936 3080 4169 3108
rect 3936 3068 3942 3080
rect 4157 3077 4169 3080
rect 4203 3077 4215 3111
rect 4157 3071 4215 3077
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 4172 3040 4200 3071
rect 4522 3068 4528 3120
rect 4580 3108 4586 3120
rect 4678 3111 4736 3117
rect 4678 3108 4690 3111
rect 4580 3080 4690 3108
rect 4580 3068 4586 3080
rect 4678 3077 4690 3080
rect 4724 3077 4736 3111
rect 6914 3108 6920 3120
rect 4678 3071 4736 3077
rect 6380 3080 6920 3108
rect 6380 3049 6408 3080
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 7466 3108 7472 3120
rect 7024 3080 7472 3108
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4172 3012 4445 3040
rect 2317 3003 2375 3009
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6632 3043 6690 3049
rect 6632 3009 6644 3043
rect 6678 3040 6690 3043
rect 7024 3040 7052 3080
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 7852 3117 7880 3148
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8996 3148 9137 3176
rect 8996 3136 9002 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9125 3139 9183 3145
rect 10229 3179 10287 3185
rect 10229 3145 10241 3179
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 7837 3111 7895 3117
rect 7837 3077 7849 3111
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 9769 3111 9827 3117
rect 9769 3077 9781 3111
rect 9815 3108 9827 3111
rect 10244 3108 10272 3139
rect 9815 3080 10272 3108
rect 9815 3077 9827 3080
rect 9769 3071 9827 3077
rect 6678 3012 7052 3040
rect 6678 3009 6690 3012
rect 6632 3003 6690 3009
rect 2332 2972 2360 3003
rect 4154 2972 4160 2984
rect 2332 2944 4160 2972
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 2406 2864 2412 2916
rect 2464 2864 2470 2916
rect 6012 2904 6040 3003
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7248 3012 10364 3040
rect 7248 3000 7254 3012
rect 8110 2932 8116 2984
rect 8168 2932 8174 2984
rect 10336 2972 10364 3012
rect 10410 3000 10416 3052
rect 10468 3000 10474 3052
rect 10502 2972 10508 2984
rect 10336 2944 10508 2972
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 7745 2907 7803 2913
rect 5368 2876 5948 2904
rect 6012 2876 6408 2904
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 5368 2836 5396 2876
rect 2924 2808 5396 2836
rect 2924 2796 2930 2808
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5813 2839 5871 2845
rect 5813 2836 5825 2839
rect 5500 2808 5825 2836
rect 5500 2796 5506 2808
rect 5813 2805 5825 2808
rect 5859 2805 5871 2839
rect 5920 2836 5948 2876
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5920 2808 6193 2836
rect 5813 2799 5871 2805
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6380 2836 6408 2876
rect 7745 2873 7757 2907
rect 7791 2904 7803 2907
rect 8128 2904 8156 2932
rect 7791 2876 8156 2904
rect 7791 2873 7803 2876
rect 7745 2867 7803 2873
rect 7466 2836 7472 2848
rect 6380 2808 7472 2836
rect 6181 2799 6239 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 7892 2808 9873 2836
rect 7892 2796 7898 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 1728 2604 2912 2632
rect 1728 2592 1734 2604
rect 1504 2536 2360 2564
rect 1504 2508 1532 2536
rect 1486 2456 1492 2508
rect 1544 2456 1550 2508
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2332 2505 2360 2536
rect 2590 2524 2596 2576
rect 2648 2524 2654 2576
rect 2133 2499 2191 2505
rect 2133 2496 2145 2499
rect 2004 2468 2145 2496
rect 2004 2456 2010 2468
rect 2133 2465 2145 2468
rect 2179 2465 2191 2499
rect 2133 2459 2191 2465
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2465 2375 2499
rect 2884 2496 2912 2604
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 6420 2604 7236 2632
rect 6420 2592 6426 2604
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 3007 2536 6914 2564
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 3881 2499 3939 2505
rect 2884 2468 3372 2496
rect 2317 2459 2375 2465
rect 1854 2428 1860 2440
rect 1688 2400 1860 2428
rect 1688 2369 1716 2400
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2866 2388 2872 2440
rect 2924 2388 2930 2440
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 3344 2428 3372 2468
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4430 2496 4436 2508
rect 3927 2468 4436 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 6886 2496 6914 2536
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6886 2468 7113 2496
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3344 2400 4261 2428
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 1673 2363 1731 2369
rect 1673 2329 1685 2363
rect 1719 2329 1731 2363
rect 1673 2323 1731 2329
rect 2038 2320 2044 2372
rect 2096 2320 2102 2372
rect 5534 2320 5540 2372
rect 5592 2320 5598 2372
rect 5629 2363 5687 2369
rect 5629 2329 5641 2363
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4341 2295 4399 2301
rect 4341 2292 4353 2295
rect 4120 2264 4353 2292
rect 4120 2252 4126 2264
rect 4341 2261 4353 2264
rect 4387 2261 4399 2295
rect 4341 2255 4399 2261
rect 5074 2252 5080 2304
rect 5132 2252 5138 2304
rect 5644 2292 5672 2323
rect 6822 2320 6828 2372
rect 6880 2360 6886 2372
rect 7208 2360 7236 2604
rect 7300 2604 8585 2632
rect 7300 2505 7328 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 7745 2567 7803 2573
rect 7745 2533 7757 2567
rect 7791 2564 7803 2567
rect 8205 2567 8263 2573
rect 8205 2564 8217 2567
rect 7791 2536 8217 2564
rect 7791 2533 7803 2536
rect 7745 2527 7803 2533
rect 8205 2533 8217 2536
rect 8251 2564 8263 2567
rect 9585 2567 9643 2573
rect 8251 2536 9076 2564
rect 8251 2533 8263 2536
rect 8205 2527 8263 2533
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7616 2468 7849 2496
rect 7616 2456 7622 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 9048 2505 9076 2536
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 10226 2564 10232 2576
rect 9631 2536 10232 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7984 2468 8033 2496
rect 7984 2456 7990 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9306 2456 9312 2508
rect 9364 2496 9370 2508
rect 9364 2468 10364 2496
rect 9364 2456 9370 2468
rect 10336 2437 10364 2468
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 10321 2431 10379 2437
rect 8757 2391 8815 2397
rect 9692 2400 9996 2428
rect 8772 2360 8800 2391
rect 6880 2332 7144 2360
rect 7208 2332 8800 2360
rect 6880 2320 6886 2332
rect 6546 2292 6552 2304
rect 5644 2264 6552 2292
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 6914 2252 6920 2304
rect 6972 2252 6978 2304
rect 7116 2292 7144 2332
rect 9122 2320 9128 2372
rect 9180 2320 9186 2372
rect 9692 2360 9720 2400
rect 9232 2332 9720 2360
rect 9232 2292 9260 2332
rect 9858 2320 9864 2372
rect 9916 2320 9922 2372
rect 9968 2360 9996 2400
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 9968 2332 10548 2360
rect 7116 2264 9260 2292
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 10520 2301 10548 2332
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9640 2264 9965 2292
rect 9640 2252 9646 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 2774 2048 2780 2100
rect 2832 2088 2838 2100
rect 9122 2088 9128 2100
rect 2832 2060 9128 2088
rect 2832 2048 2838 2060
rect 9122 2048 9128 2060
rect 9180 2048 9186 2100
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 6552 9664 6604 9716
rect 1768 9596 1820 9648
rect 2964 9596 3016 9648
rect 4160 9596 4212 9648
rect 940 9528 992 9580
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 2688 9460 2740 9512
rect 2964 9460 3016 9512
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 5724 9528 5776 9580
rect 9588 9664 9640 9716
rect 8944 9596 8996 9648
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 1400 9367 1452 9376
rect 1400 9333 1409 9367
rect 1409 9333 1443 9367
rect 1443 9333 1452 9367
rect 1400 9324 1452 9333
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 5356 9392 5408 9444
rect 7748 9392 7800 9444
rect 9220 9460 9272 9512
rect 10508 9528 10560 9580
rect 10048 9392 10100 9444
rect 10140 9392 10192 9444
rect 7840 9324 7892 9376
rect 9036 9324 9088 9376
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 572 9120 624 9172
rect 1952 9120 2004 9172
rect 2688 9120 2740 9172
rect 4344 9120 4396 9172
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 9312 9120 9364 9172
rect 9956 9052 10008 9104
rect 1492 8891 1544 8900
rect 1492 8857 1501 8891
rect 1501 8857 1535 8891
rect 1535 8857 1544 8891
rect 1492 8848 1544 8857
rect 4252 8916 4304 8968
rect 9588 8891 9640 8900
rect 9588 8857 9597 8891
rect 9597 8857 9631 8891
rect 9631 8857 9640 8891
rect 9588 8848 9640 8857
rect 11336 8916 11388 8968
rect 10140 8891 10192 8900
rect 10140 8857 10149 8891
rect 10149 8857 10183 8891
rect 10183 8857 10192 8891
rect 10140 8848 10192 8857
rect 2044 8780 2096 8832
rect 6644 8780 6696 8832
rect 9220 8780 9272 8832
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 1400 8576 1452 8628
rect 2044 8576 2096 8628
rect 9128 8576 9180 8628
rect 9588 8576 9640 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 9404 8508 9456 8560
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 1768 8304 1820 8356
rect 7472 8372 7524 8424
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 6920 8304 6972 8356
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 9956 8372 10008 8424
rect 9220 8236 9272 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 5540 8032 5592 8084
rect 5632 8032 5684 8084
rect 6276 7896 6328 7948
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 9404 7896 9456 7948
rect 9956 7828 10008 7880
rect 9864 7760 9916 7812
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 5356 7692 5408 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 6828 7692 6880 7744
rect 7840 7692 7892 7744
rect 8116 7692 8168 7744
rect 8668 7692 8720 7744
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 5172 7488 5224 7540
rect 6368 7488 6420 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 1492 7284 1544 7336
rect 5356 7352 5408 7404
rect 8668 7488 8720 7540
rect 9956 7488 10008 7540
rect 9312 7420 9364 7472
rect 6828 7352 6880 7404
rect 7656 7352 7708 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9220 7352 9272 7404
rect 9404 7352 9456 7404
rect 10876 7352 10928 7404
rect 2504 7216 2556 7268
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 7656 7216 7708 7268
rect 7840 7216 7892 7268
rect 2872 7148 2924 7200
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 8668 7148 8720 7200
rect 8852 7148 8904 7200
rect 10048 7216 10100 7268
rect 10416 7148 10468 7200
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 2320 6944 2372 6996
rect 2504 6876 2556 6928
rect 1860 6740 1912 6792
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 6460 6919 6512 6928
rect 6460 6885 6469 6919
rect 6469 6885 6503 6919
rect 6503 6885 6512 6919
rect 6460 6876 6512 6885
rect 3884 6808 3936 6860
rect 7380 6944 7432 6996
rect 7656 6876 7708 6928
rect 9220 6944 9272 6996
rect 6828 6808 6880 6860
rect 7288 6808 7340 6860
rect 3240 6672 3292 6724
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 1952 6604 2004 6656
rect 2504 6604 2556 6656
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3700 6604 3752 6656
rect 5816 6740 5868 6792
rect 6276 6740 6328 6792
rect 6368 6672 6420 6724
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9036 6740 9088 6792
rect 6184 6604 6236 6656
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 7564 6604 7616 6656
rect 9404 6672 9456 6724
rect 9680 6604 9732 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 1768 6332 1820 6384
rect 2320 6400 2372 6452
rect 2412 6400 2464 6452
rect 3056 6400 3108 6452
rect 3148 6400 3200 6452
rect 940 6264 992 6316
rect 2412 6196 2464 6248
rect 1676 6171 1728 6180
rect 1676 6137 1685 6171
rect 1685 6137 1719 6171
rect 1719 6137 1728 6171
rect 1676 6128 1728 6137
rect 1584 6060 1636 6112
rect 5172 6400 5224 6452
rect 5724 6400 5776 6452
rect 6552 6400 6604 6452
rect 7748 6400 7800 6452
rect 8944 6400 8996 6452
rect 4988 6332 5040 6384
rect 5540 6332 5592 6384
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 3884 6264 3936 6316
rect 6092 6332 6144 6384
rect 6276 6332 6328 6384
rect 6460 6332 6512 6384
rect 7288 6264 7340 6316
rect 8668 6264 8720 6316
rect 6276 6196 6328 6248
rect 6368 6196 6420 6248
rect 7564 6196 7616 6248
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10324 6264 10376 6316
rect 3148 6128 3200 6180
rect 3516 6128 3568 6180
rect 3240 6060 3292 6112
rect 3700 6060 3752 6112
rect 4436 6060 4488 6112
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 9404 6128 9456 6180
rect 7840 6060 7892 6112
rect 9220 6060 9272 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 10232 6060 10284 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1860 5856 1912 5908
rect 2780 5856 2832 5908
rect 4436 5856 4488 5908
rect 5080 5856 5132 5908
rect 2044 5652 2096 5704
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 2780 5652 2832 5704
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 3332 5652 3384 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4068 5788 4120 5840
rect 5724 5788 5776 5840
rect 6184 5856 6236 5908
rect 6276 5856 6328 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 4344 5652 4396 5704
rect 5540 5652 5592 5704
rect 6092 5720 6144 5772
rect 7840 5788 7892 5840
rect 6736 5720 6788 5772
rect 6828 5652 6880 5704
rect 6920 5652 6972 5704
rect 8852 5856 8904 5908
rect 10048 5856 10100 5908
rect 9128 5720 9180 5772
rect 9956 5788 10008 5840
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 2044 5516 2096 5568
rect 2688 5516 2740 5568
rect 6184 5584 6236 5636
rect 2872 5516 2924 5568
rect 3700 5516 3752 5568
rect 4160 5516 4212 5568
rect 4712 5516 4764 5568
rect 5632 5516 5684 5568
rect 8116 5584 8168 5636
rect 7380 5516 7432 5568
rect 8392 5584 8444 5636
rect 9956 5584 10008 5636
rect 9404 5516 9456 5568
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 1768 5312 1820 5364
rect 940 5176 992 5228
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2872 5244 2924 5296
rect 3148 5244 3200 5296
rect 3056 5108 3108 5160
rect 3792 5312 3844 5364
rect 4712 5312 4764 5364
rect 4896 5312 4948 5364
rect 4252 5176 4304 5228
rect 4344 5176 4396 5228
rect 5080 5312 5132 5364
rect 6092 5312 6144 5364
rect 8760 5312 8812 5364
rect 5356 5176 5408 5228
rect 5632 5176 5684 5228
rect 6736 5176 6788 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8668 5219 8720 5228
rect 8668 5185 8702 5219
rect 8702 5185 8720 5219
rect 8668 5176 8720 5185
rect 8944 5176 8996 5228
rect 3148 5040 3200 5092
rect 1768 4972 1820 5024
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6920 5040 6972 5092
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 10140 4972 10192 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 2780 4768 2832 4820
rect 3148 4768 3200 4820
rect 3700 4768 3752 4820
rect 1952 4632 2004 4684
rect 2872 4632 2924 4684
rect 5540 4743 5592 4752
rect 5540 4709 5549 4743
rect 5549 4709 5583 4743
rect 5583 4709 5592 4743
rect 5540 4700 5592 4709
rect 6092 4700 6144 4752
rect 6920 4743 6972 4752
rect 6920 4709 6929 4743
rect 6929 4709 6963 4743
rect 6963 4709 6972 4743
rect 6920 4700 6972 4709
rect 2044 4564 2096 4616
rect 2228 4564 2280 4616
rect 3056 4564 3108 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4344 4564 4396 4616
rect 4620 4564 4672 4616
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5448 4564 5500 4616
rect 5724 4564 5776 4616
rect 8392 4632 8444 4684
rect 8668 4768 8720 4820
rect 9404 4700 9456 4752
rect 9128 4632 9180 4684
rect 9956 4700 10008 4752
rect 10048 4632 10100 4684
rect 1308 4428 1360 4480
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 3148 4428 3200 4480
rect 4344 4428 4396 4480
rect 4528 4428 4580 4480
rect 6828 4496 6880 4548
rect 6920 4496 6972 4548
rect 8668 4496 8720 4548
rect 7380 4428 7432 4480
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1952 4267 2004 4276
rect 1952 4233 1961 4267
rect 1961 4233 1995 4267
rect 1995 4233 2004 4267
rect 1952 4224 2004 4233
rect 2136 4224 2188 4276
rect 3792 4224 3844 4276
rect 4068 4224 4120 4276
rect 2412 4088 2464 4140
rect 4620 4224 4672 4276
rect 5080 4224 5132 4276
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4804 4088 4856 4140
rect 5540 4088 5592 4140
rect 6828 4156 6880 4208
rect 7472 4156 7524 4208
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 10048 4224 10100 4276
rect 9956 4156 10008 4208
rect 8116 4088 8168 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 1676 3952 1728 4004
rect 1952 3952 2004 4004
rect 388 3884 440 3936
rect 4896 4020 4948 4072
rect 3976 3952 4028 4004
rect 5264 4020 5316 4072
rect 7472 4020 7524 4072
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 9956 4020 10008 4072
rect 6276 3952 6328 4004
rect 3884 3884 3936 3936
rect 4344 3884 4396 3936
rect 4804 3884 4856 3936
rect 4988 3884 5040 3936
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5632 3884 5684 3936
rect 6368 3884 6420 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 7932 3884 7984 3936
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 2044 3680 2096 3732
rect 2596 3544 2648 3596
rect 3056 3680 3108 3732
rect 4160 3680 4212 3732
rect 4436 3680 4488 3732
rect 4620 3680 4672 3732
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 5540 3680 5592 3732
rect 6920 3680 6972 3732
rect 7932 3680 7984 3732
rect 8024 3680 8076 3732
rect 2780 3612 2832 3664
rect 5448 3612 5500 3664
rect 6184 3612 6236 3664
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 2412 3451 2464 3460
rect 2412 3417 2421 3451
rect 2421 3417 2455 3451
rect 2455 3417 2464 3451
rect 2412 3408 2464 3417
rect 3516 3408 3568 3460
rect 4344 3476 4396 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5080 3476 5132 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 10324 3655 10376 3664
rect 10324 3621 10333 3655
rect 10333 3621 10367 3655
rect 10367 3621 10376 3655
rect 10324 3612 10376 3621
rect 1584 3340 1636 3392
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 5448 3340 5500 3392
rect 5724 3408 5776 3460
rect 7196 3340 7248 3392
rect 7288 3340 7340 3392
rect 9864 3451 9916 3460
rect 9864 3417 9873 3451
rect 9873 3417 9907 3451
rect 9907 3417 9916 3451
rect 9864 3408 9916 3417
rect 9036 3340 9088 3392
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 1400 3136 1452 3188
rect 2504 3136 2556 3188
rect 7656 3136 7708 3188
rect 3884 3068 3936 3120
rect 4528 3068 4580 3120
rect 6920 3068 6972 3120
rect 7472 3068 7524 3120
rect 8944 3136 8996 3188
rect 4160 2932 4212 2984
rect 2412 2907 2464 2916
rect 2412 2873 2421 2907
rect 2421 2873 2455 2907
rect 2455 2873 2464 2907
rect 2412 2864 2464 2873
rect 7196 3000 7248 3052
rect 8116 2932 8168 2984
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 10508 2932 10560 2984
rect 2872 2796 2924 2848
rect 5448 2796 5500 2848
rect 7472 2796 7524 2848
rect 7840 2796 7892 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 1676 2592 1728 2644
rect 1492 2456 1544 2508
rect 1952 2456 2004 2508
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 6368 2592 6420 2644
rect 1860 2388 1912 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4436 2456 4488 2508
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 5172 2388 5224 2440
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 4068 2252 4120 2304
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 6828 2320 6880 2372
rect 7564 2456 7616 2508
rect 7932 2456 7984 2508
rect 10232 2524 10284 2576
rect 9312 2456 9364 2508
rect 6552 2252 6604 2304
rect 6920 2295 6972 2304
rect 6920 2261 6929 2295
rect 6929 2261 6963 2295
rect 6963 2261 6972 2295
rect 6920 2252 6972 2261
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 9864 2363 9916 2372
rect 9864 2329 9873 2363
rect 9873 2329 9907 2363
rect 9907 2329 9916 2363
rect 9864 2320 9916 2329
rect 9588 2252 9640 2304
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 2780 2048 2832 2100
rect 9128 2048 9180 2100
<< metal2 >>
rect 570 11200 626 12000
rect 1766 11200 1822 12000
rect 2962 11200 3018 12000
rect 4158 11200 4214 12000
rect 5354 11200 5410 12000
rect 6550 11200 6606 12000
rect 7746 11200 7802 12000
rect 8942 11200 8998 12000
rect 9310 11248 9366 11257
rect 584 9178 612 11200
rect 1780 9654 1808 11200
rect 2778 10160 2834 10169
rect 2778 10095 2834 10104
rect 2792 9674 2820 10095
rect 1768 9648 1820 9654
rect 2700 9646 2820 9674
rect 2976 9654 3004 11200
rect 3054 10976 3110 10985
rect 3054 10911 3110 10920
rect 2964 9648 3016 9654
rect 1768 9590 1820 9596
rect 2410 9616 2466 9625
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 1952 9580 2004 9586
rect 2410 9551 2412 9560
rect 1952 9522 2004 9528
rect 2464 9551 2466 9560
rect 2412 9522 2464 9528
rect 572 9172 624 9178
rect 572 9114 624 9120
rect 952 9081 980 9522
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1412 8634 1440 9318
rect 1964 9178 1992 9522
rect 2700 9518 2728 9646
rect 3068 9625 3096 10911
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 4172 9654 4200 11200
rect 4160 9648 4212 9654
rect 2964 9590 3016 9596
rect 3054 9616 3110 9625
rect 4160 9590 4212 9596
rect 3054 9551 3110 9560
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 2688 9512 2740 9518
rect 2964 9512 3016 9518
rect 2688 9454 2740 9460
rect 2792 9472 2964 9500
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 2700 9178 2728 9318
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1504 8401 1532 8842
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8634 2084 8774
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1490 8392 1546 8401
rect 1490 8327 1546 8336
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1504 6474 1532 7278
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1412 6446 1532 6474
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 5817 980 6258
rect 938 5808 994 5817
rect 938 5743 994 5752
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4729 980 5170
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1308 4480 1360 4486
rect 1308 4422 1360 4428
rect 388 3936 440 3942
rect 388 3878 440 3884
rect 400 800 428 3878
rect 1320 800 1348 4422
rect 1412 3194 1440 6446
rect 1688 6304 1716 6598
rect 1780 6390 1808 8298
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 6798 1900 7346
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1504 6276 1716 6304
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1504 2514 1532 6276
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 3482 1624 6054
rect 1688 5681 1716 6122
rect 1674 5672 1730 5681
rect 1674 5607 1730 5616
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1688 4010 1716 5510
rect 1780 5370 1808 6326
rect 1872 5914 1900 6734
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1964 5273 1992 6598
rect 2056 5710 2084 8570
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2332 6458 2360 6938
rect 2516 6934 2544 7210
rect 2504 6928 2556 6934
rect 2792 6882 2820 9472
rect 2964 9454 3016 9460
rect 4356 9178 4384 9522
rect 5368 9450 5396 11200
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 6564 9722 6592 11200
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2504 6870 2556 6876
rect 2516 6746 2544 6870
rect 2424 6718 2544 6746
rect 2700 6854 2820 6882
rect 2424 6458 2452 6718
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2424 6254 2452 6287
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 1950 5264 2006 5273
rect 1860 5228 1912 5234
rect 1950 5199 2006 5208
rect 1860 5170 1912 5176
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1780 3890 1808 4966
rect 1872 4162 1900 5170
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1964 4282 1992 4626
rect 2056 4622 2084 5510
rect 2332 5137 2360 5646
rect 2318 5128 2374 5137
rect 2318 5063 2374 5072
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4282 2176 4422
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2240 4162 2268 4558
rect 2516 4162 2544 6598
rect 1872 4134 2268 4162
rect 2424 4146 2544 4162
rect 2412 4140 2544 4146
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1780 3862 1900 3890
rect 1596 3454 1716 3482
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 2553 1624 3334
rect 1688 2650 1716 3454
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1582 2544 1638 2553
rect 1492 2508 1544 2514
rect 1582 2479 1638 2488
rect 1492 2450 1544 2456
rect 1872 2446 1900 3862
rect 1964 2514 1992 3946
rect 2056 3738 2084 4134
rect 2464 4134 2544 4140
rect 2608 4162 2636 6598
rect 2700 5574 2728 6854
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 5914 2820 6734
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 5710 2912 7142
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3056 6792 3108 6798
rect 3054 6760 3056 6769
rect 3108 6760 3110 6769
rect 3054 6695 3110 6704
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 2976 6582 3188 6610
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2792 5114 2820 5646
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5302 2912 5510
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2792 5086 2912 5114
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4826 2820 4966
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2884 4690 2912 5086
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2870 4584 2926 4593
rect 2870 4519 2926 4528
rect 2608 4134 2820 4162
rect 2412 4082 2464 4088
rect 2502 4040 2558 4049
rect 2502 3975 2558 3984
rect 2686 4040 2742 4049
rect 2686 3975 2742 3984
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2410 3496 2466 3505
rect 2410 3431 2412 3440
rect 2464 3431 2466 3440
rect 2412 3402 2464 3408
rect 2516 3194 2544 3975
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2410 2952 2466 2961
rect 2410 2887 2412 2896
rect 2464 2887 2466 2896
rect 2412 2858 2464 2864
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2608 2582 2636 3538
rect 2700 3534 2728 3975
rect 2792 3670 2820 4134
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 2056 1170 2084 2314
rect 2792 2106 2820 3334
rect 2884 2854 2912 4519
rect 2976 3641 3004 6582
rect 3160 6458 3188 6582
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3068 5409 3096 6394
rect 3252 6202 3280 6666
rect 3700 6656 3752 6662
rect 3752 6616 3832 6644
rect 3700 6598 3752 6604
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3148 6180 3200 6186
rect 3252 6174 3372 6202
rect 3148 6122 3200 6128
rect 3054 5400 3110 5409
rect 3054 5335 3110 5344
rect 3160 5302 3188 6122
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5953 3280 6054
rect 3238 5944 3294 5953
rect 3238 5879 3294 5888
rect 3344 5710 3372 6174
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3528 5817 3556 6122
rect 3514 5808 3570 5817
rect 3514 5743 3570 5752
rect 3332 5704 3384 5710
rect 3238 5672 3294 5681
rect 3620 5681 3648 6258
rect 3804 6225 3832 6616
rect 3896 6322 3924 6802
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3332 5646 3384 5652
rect 3606 5672 3662 5681
rect 3238 5607 3294 5616
rect 3606 5607 3662 5616
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4706 3096 5102
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3160 4826 3188 5034
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3068 4678 3188 4706
rect 3056 4616 3108 4622
rect 3054 4584 3056 4593
rect 3108 4584 3110 4593
rect 3054 4519 3110 4528
rect 3160 4486 3188 4678
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3068 3738 3096 4422
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2962 3632 3018 3641
rect 2962 3567 3018 3576
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2446 2912 2790
rect 3252 2446 3280 5607
rect 3712 5574 3740 6054
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3804 5370 3832 5646
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4826 3740 5102
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3804 4282 3832 4558
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3896 3942 3924 6258
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 3988 4010 4016 4927
rect 4080 4282 4108 5782
rect 4172 5574 4200 5879
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4264 5352 4292 8910
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 5552 8090 5580 9522
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5184 7546 5212 7686
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5368 7410 5396 7686
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4436 6112 4488 6118
rect 4356 6072 4436 6100
rect 4356 5710 4384 6072
rect 4436 6054 4488 6060
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4172 5324 4292 5352
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3936 3936 3942
rect 3514 3904 3570 3913
rect 3884 3878 3936 3884
rect 3514 3839 3570 3848
rect 3528 3466 3556 3839
rect 3516 3460 3568 3466
rect 3516 3402 3568 3408
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3896 3126 3924 3878
rect 4172 3738 4200 5324
rect 4356 5234 4384 5646
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4264 4146 4292 5170
rect 4356 4622 4384 5170
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4321 4384 4422
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4448 4196 4476 5850
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5370 4752 5510
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4896 5364 4948 5370
rect 5000 5352 5028 6326
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5092 5370 5120 5850
rect 4948 5324 5028 5352
rect 5080 5364 5132 5370
rect 4896 5306 4948 5312
rect 5080 5306 5132 5312
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4356 4168 4476 4196
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4356 4060 4384 4168
rect 4356 4032 4476 4060
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 4172 2990 4200 3674
rect 4356 3534 4384 3878
rect 4448 3738 4476 4032
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4448 2514 4476 3470
rect 4540 3126 4568 4422
rect 4632 4282 4660 4558
rect 4802 4312 4858 4321
rect 4620 4276 4672 4282
rect 4858 4270 4936 4298
rect 5092 4282 5120 4558
rect 4802 4247 4858 4256
rect 4620 4218 4672 4224
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3942 4844 4082
rect 4908 4078 4936 4270
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 5000 3738 5028 3878
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4632 3534 4660 3674
rect 5078 3632 5134 3641
rect 5078 3567 5134 3576
rect 5092 3534 5120 3567
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 5184 2446 5212 6394
rect 5540 6384 5592 6390
rect 5262 6352 5318 6361
rect 5644 6372 5672 8026
rect 5736 6458 5764 9522
rect 7760 9450 7788 11200
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 8956 9654 8984 11200
rect 10138 11200 10194 12000
rect 11334 11200 11390 12000
rect 9310 11183 9366 11192
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6798 5856 7142
rect 6288 6798 6316 7890
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7546 6408 7686
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5592 6344 5672 6372
rect 6092 6384 6144 6390
rect 5540 6326 5592 6332
rect 6092 6326 6144 6332
rect 5262 6287 5318 6296
rect 5276 4078 5304 6287
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5953 5856 6054
rect 5814 5944 5870 5953
rect 5814 5879 5870 5888
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5250 5580 5646
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5368 5234 5580 5250
rect 5644 5234 5672 5510
rect 5356 5228 5580 5234
rect 5408 5222 5580 5228
rect 5632 5228 5684 5234
rect 5356 5170 5408 5176
rect 5632 5170 5684 5176
rect 5540 5160 5592 5166
rect 5460 5108 5540 5114
rect 5460 5102 5592 5108
rect 5630 5128 5686 5137
rect 5460 5086 5580 5102
rect 5460 4622 5488 5086
rect 5630 5063 5686 5072
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5552 4146 5580 4694
rect 5644 4434 5672 5063
rect 5736 4622 5764 5782
rect 6104 5778 6132 6326
rect 6196 5914 6224 6598
rect 6288 6390 6316 6734
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6380 6254 6408 6666
rect 6472 6390 6500 6870
rect 6564 6458 6592 7822
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6550 6216 6606 6225
rect 6288 5914 6316 6190
rect 6550 6151 6606 6160
rect 6564 5930 6592 6151
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6380 5902 6592 5930
rect 6274 5808 6330 5817
rect 6092 5772 6144 5778
rect 6274 5743 6330 5752
rect 6092 5714 6144 5720
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6104 4758 6132 5306
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5644 4406 5764 4434
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5264 4072 5316 4078
rect 5316 4032 5396 4060
rect 5264 4014 5316 4020
rect 5368 3534 5396 4032
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5460 3670 5488 3878
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 2836 5396 3470
rect 5460 3398 5488 3606
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5448 2848 5500 2854
rect 5368 2808 5448 2836
rect 5448 2790 5500 2796
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5552 2378 5580 3674
rect 5644 3097 5672 3878
rect 5736 3466 5764 4406
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 6196 3670 6224 5578
rect 6288 4729 6316 5743
rect 6274 4720 6330 4729
rect 6380 4706 6408 5902
rect 6380 4678 6592 4706
rect 6274 4655 6330 4664
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 5630 3088 5686 3097
rect 5630 3023 5686 3032
rect 6196 2514 6224 3606
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 3332 2304 3384 2310
rect 3160 2264 3332 2292
rect 2780 2100 2832 2106
rect 2780 2042 2832 2048
rect 2056 1142 2268 1170
rect 2240 800 2268 1142
rect 3160 800 3188 2264
rect 4068 2304 4120 2310
rect 3332 2246 3384 2252
rect 3988 2264 4068 2292
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3988 1170 4016 2264
rect 5080 2304 5132 2310
rect 4068 2246 4120 2252
rect 5000 2264 5080 2292
rect 3988 1142 4108 1170
rect 4080 800 4108 1142
rect 5000 800 5028 2264
rect 5080 2246 5132 2252
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 5920 870 6040 898
rect 5920 800 5948 870
rect 386 0 442 800
rect 1306 0 1362 800
rect 2226 0 2282 800
rect 3146 0 3202 800
rect 4066 0 4122 800
rect 4986 0 5042 800
rect 5906 0 5962 800
rect 6012 762 6040 870
rect 6288 762 6316 3946
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 2650 6408 3878
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6564 2310 6592 4678
rect 6656 2446 6684 8774
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 7410 6868 7686
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 6866 6868 7346
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6734 5944 6790 5953
rect 6734 5879 6790 5888
rect 6748 5778 6776 5879
rect 6932 5794 6960 8298
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7392 7002 7420 7822
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6860 7340 6866
rect 7340 6820 7420 6848
rect 7288 6802 7340 6808
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6322 7328 6598
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6840 5766 6960 5794
rect 6840 5710 6868 5766
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6748 1465 6776 5170
rect 6932 5098 6960 5646
rect 7392 5574 7420 6820
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6932 4758 6960 5034
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6840 4214 6868 4490
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6840 2378 6868 4150
rect 6932 3738 6960 4490
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6932 3126 6960 3674
rect 7286 3496 7342 3505
rect 7286 3431 7342 3440
rect 7300 3398 7328 3431
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7208 3058 7236 3334
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7392 2938 7420 4422
rect 7484 4214 7512 8366
rect 7668 7410 7696 8366
rect 7852 7750 7880 9318
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 6934 7696 7210
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6254 7604 6598
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7668 5914 7696 6870
rect 7760 6458 7788 7278
rect 7852 7274 7880 7686
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7852 5846 7880 6054
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 8128 5794 8156 7686
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8680 7546 8708 7686
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8680 6322 8708 7142
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8206 5808 8262 5817
rect 8128 5766 8206 5794
rect 8206 5743 8262 5752
rect 8772 5658 8800 8434
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 5914 8892 7142
rect 9048 6798 9076 9318
rect 9140 8634 9168 9522
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9178 9260 9454
rect 9324 9178 9352 11183
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9600 9722 9628 10095
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 10152 9450 10180 11200
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9968 9110 9996 9318
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9232 8498 9260 8774
rect 9600 8634 9628 8842
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9404 8560 9456 8566
rect 9968 8514 9996 9046
rect 9404 8502 9456 8508
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7410 9260 8230
rect 9416 7954 9444 8502
rect 9876 8498 9996 8514
rect 9864 8492 9996 8498
rect 9916 8486 9996 8492
rect 9864 8434 9916 8440
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9968 7993 9996 8366
rect 9954 7984 10010 7993
rect 9404 7948 9456 7954
rect 9954 7919 10010 7928
rect 9404 7890 9456 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 8956 6458 8984 6734
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8116 5636 8168 5642
rect 8392 5636 8444 5642
rect 8168 5596 8392 5624
rect 8116 5578 8168 5584
rect 8772 5630 8892 5658
rect 8392 5578 8444 5584
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3126 7512 4014
rect 7668 3194 7696 4966
rect 8404 4690 8432 5170
rect 8680 4826 8708 5170
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8680 4282 8708 4490
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 4072 8076 4078
rect 8022 4040 8024 4049
rect 8076 4040 8078 4049
rect 8022 3975 8078 3984
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7760 3346 7788 3878
rect 7944 3738 7972 3878
rect 8036 3738 8064 3975
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7760 3318 7972 3346
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7392 2910 7604 2938
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7484 2553 7512 2790
rect 7470 2544 7526 2553
rect 7576 2514 7604 2910
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7470 2479 7526 2488
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6734 1456 6790 1465
rect 6932 1442 6960 2246
rect 7852 1442 7880 2790
rect 7944 2514 7972 3318
rect 8128 2990 8156 4082
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8772 2530 8800 5306
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8680 2502 8800 2530
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 6734 1391 6790 1400
rect 6840 1414 6960 1442
rect 7760 1414 7880 1442
rect 6840 800 6868 1414
rect 7760 800 7788 1414
rect 8680 800 8708 2502
rect 8864 1442 8892 5630
rect 8956 5234 8984 6394
rect 9140 5778 9168 7346
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9324 6458 9352 7414
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 6730 9444 7346
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9232 6118 9260 6258
rect 9416 6186 9444 6666
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9876 6202 9904 7754
rect 9968 7546 9996 7822
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 10060 7274 10088 9386
rect 10520 9081 10548 9522
rect 10506 9072 10562 9081
rect 10506 9007 10562 9016
rect 11348 8974 11376 11200
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9404 6180 9456 6186
rect 9876 6174 9996 6202
rect 9404 6122 9456 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9034 5264 9090 5273
rect 8944 5228 8996 5234
rect 9034 5199 9090 5208
rect 8944 5170 8996 5176
rect 8956 3194 8984 5170
rect 9048 3398 9076 5199
rect 9140 4690 9168 5714
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 4758 9444 5510
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9678 4720 9734 4729
rect 9128 4684 9180 4690
rect 9734 4678 9812 4706
rect 9678 4655 9734 4664
rect 9128 4626 9180 4632
rect 9784 4026 9812 4678
rect 9876 4146 9904 6054
rect 9968 5846 9996 6174
rect 10060 5914 10088 6258
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9968 4758 9996 5578
rect 10152 5030 10180 8842
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9968 4214 9996 4694
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4282 10088 4626
rect 10152 4593 10180 4966
rect 10138 4584 10194 4593
rect 10138 4519 10194 4528
rect 10244 4434 10272 6054
rect 10152 4406 10272 4434
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9956 4072 10008 4078
rect 9784 3998 9904 4026
rect 9956 4014 10008 4020
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9876 3466 9904 3998
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9968 2961 9996 4014
rect 9954 2952 10010 2961
rect 9954 2887 10010 2896
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9140 2106 9168 2314
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 8942 1456 8998 1465
rect 8864 1414 8942 1442
rect 8942 1391 8998 1400
rect 6012 734 6316 762
rect 6826 0 6882 800
rect 7746 0 7802 800
rect 8666 0 8722 800
rect 9324 377 9352 2450
rect 9864 2372 9916 2378
rect 10152 2360 10180 4406
rect 10336 3670 10364 6258
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10336 2774 10364 3606
rect 10428 3058 10456 7142
rect 10888 6905 10916 7346
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10244 2746 10364 2774
rect 10244 2582 10272 2746
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 9916 2332 10180 2360
rect 9864 2314 9916 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9600 800 9628 2246
rect 10520 800 10548 2926
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 9310 368 9366 377
rect 9310 303 9366 312
rect 9586 0 9642 800
rect 10506 0 10562 800
<< via2 >>
rect 2778 10104 2834 10160
rect 3054 10920 3110 10976
rect 2410 9580 2466 9616
rect 2410 9560 2412 9580
rect 2412 9560 2464 9580
rect 2464 9560 2466 9580
rect 938 9016 994 9072
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 3054 9560 3110 9616
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 1490 8336 1546 8392
rect 1398 8200 1454 8256
rect 1398 6840 1454 6896
rect 938 5752 994 5808
rect 938 4664 994 4720
rect 1674 5616 1730 5672
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 2410 6296 2466 6352
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 1950 5208 2006 5264
rect 2318 5072 2374 5128
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 1582 2488 1638 2544
rect 3054 6740 3056 6760
rect 3056 6740 3108 6760
rect 3108 6740 3110 6760
rect 3054 6704 3110 6740
rect 2870 4528 2926 4584
rect 2502 3984 2558 4040
rect 2686 3984 2742 4040
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2410 3460 2466 3496
rect 2410 3440 2412 3460
rect 2412 3440 2464 3460
rect 2464 3440 2466 3460
rect 2410 2916 2466 2952
rect 2410 2896 2412 2916
rect 2412 2896 2464 2916
rect 2464 2896 2466 2916
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3054 5344 3110 5400
rect 3238 5888 3294 5944
rect 3514 5752 3570 5808
rect 3238 5616 3294 5672
rect 3790 6160 3846 6216
rect 3606 5616 3662 5672
rect 3054 4564 3056 4584
rect 3056 4564 3108 4584
rect 3108 4564 3110 4584
rect 3054 4528 3110 4564
rect 2962 3576 3018 3632
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 4158 5888 4214 5944
rect 3974 4936 4030 4992
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 3514 3848 3570 3904
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 4342 4256 4398 4312
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4802 4256 4858 4312
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 5078 3576 5134 3632
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 5262 6296 5318 6352
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 9310 11192 9366 11248
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 5814 5888 5870 5944
rect 5630 5072 5686 5128
rect 6550 6160 6606 6216
rect 6274 5752 6330 5808
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 6274 4664 6330 4720
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 5630 3032 5686 3088
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 6734 5888 6790 5944
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7286 3440 7342 3496
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 8206 5752 8262 5808
rect 9586 10104 9642 10160
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 9954 7928 10010 7984
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 8022 4020 8024 4040
rect 8024 4020 8076 4040
rect 8076 4020 8078 4040
rect 8022 3984 8078 4020
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 7470 2488 7526 2544
rect 6734 1400 6790 1456
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10506 9016 10562 9072
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 9034 5208 9090 5264
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 9678 4664 9734 4720
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 10138 4528 10194 4584
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9954 2896 10010 2952
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 8942 1400 8998 1456
rect 10874 6840 10930 6896
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 9310 312 9366 368
<< metal3 >>
rect 0 11250 800 11280
rect 9305 11250 9371 11253
rect 11200 11250 12000 11280
rect 0 11190 1410 11250
rect 0 11160 800 11190
rect 1350 10978 1410 11190
rect 9305 11248 12000 11250
rect 9305 11192 9310 11248
rect 9366 11192 12000 11248
rect 9305 11190 12000 11192
rect 9305 11187 9371 11190
rect 11200 11160 12000 11190
rect 3049 10978 3115 10981
rect 1350 10976 3115 10978
rect 1350 10920 3054 10976
rect 3110 10920 3115 10976
rect 1350 10918 3115 10920
rect 3049 10915 3115 10918
rect 0 10162 800 10192
rect 2773 10162 2839 10165
rect 0 10160 2839 10162
rect 0 10104 2778 10160
rect 2834 10104 2839 10160
rect 0 10102 2839 10104
rect 0 10072 800 10102
rect 2773 10099 2839 10102
rect 9581 10162 9647 10165
rect 11200 10162 12000 10192
rect 9581 10160 12000 10162
rect 9581 10104 9586 10160
rect 9642 10104 12000 10160
rect 9581 10102 12000 10104
rect 9581 10099 9647 10102
rect 11200 10072 12000 10102
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 10698 9759 11014 9760
rect 2405 9618 2471 9621
rect 3049 9618 3115 9621
rect 2405 9616 3115 9618
rect 2405 9560 2410 9616
rect 2466 9560 3054 9616
rect 3110 9560 3115 9616
rect 2405 9558 3115 9560
rect 2405 9555 2471 9558
rect 3049 9555 3115 9558
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 10501 9074 10567 9077
rect 11200 9074 12000 9104
rect 10501 9072 12000 9074
rect 10501 9016 10506 9072
rect 10562 9016 12000 9072
rect 10501 9014 12000 9016
rect 10501 9011 10567 9014
rect 11200 8984 12000 9014
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 10698 8671 11014 8672
rect 1485 8394 1551 8397
rect 1894 8394 1900 8396
rect 1485 8392 1900 8394
rect 1485 8336 1490 8392
rect 1546 8336 1900 8392
rect 1485 8334 1900 8336
rect 1485 8331 1551 8334
rect 1894 8332 1900 8334
rect 1964 8332 1970 8396
rect 1393 8258 1459 8261
rect 798 8256 1459 8258
rect 798 8200 1398 8256
rect 1454 8200 1459 8256
rect 798 8198 1459 8200
rect 798 8016 858 8198
rect 1393 8195 1459 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 9479 8127 9795 8128
rect 0 7926 858 8016
rect 9949 7986 10015 7989
rect 11200 7986 12000 8016
rect 9949 7984 12000 7986
rect 9949 7928 9954 7984
rect 10010 7928 12000 7984
rect 9949 7926 12000 7928
rect 0 7896 800 7926
rect 9949 7923 10015 7926
rect 11200 7896 12000 7926
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 10698 7583 11014 7584
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 10869 6898 10935 6901
rect 11200 6898 12000 6928
rect 10869 6896 12000 6898
rect 10869 6840 10874 6896
rect 10930 6840 12000 6896
rect 10869 6838 12000 6840
rect 10869 6835 10935 6838
rect 11200 6808 12000 6838
rect 3049 6762 3115 6765
rect 3182 6762 3188 6764
rect 3049 6760 3188 6762
rect 3049 6704 3054 6760
rect 3110 6704 3188 6760
rect 3049 6702 3188 6704
rect 3049 6699 3115 6702
rect 3182 6700 3188 6702
rect 3252 6700 3258 6764
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 10698 6495 11014 6496
rect 2405 6354 2471 6357
rect 5257 6354 5323 6357
rect 2405 6352 5323 6354
rect 2405 6296 2410 6352
rect 2466 6296 5262 6352
rect 5318 6296 5323 6352
rect 2405 6294 5323 6296
rect 2405 6291 2471 6294
rect 5257 6291 5323 6294
rect 3785 6218 3851 6221
rect 6545 6218 6611 6221
rect 3785 6216 6611 6218
rect 3785 6160 3790 6216
rect 3846 6160 6550 6216
rect 6606 6160 6611 6216
rect 3785 6158 6611 6160
rect 3785 6155 3851 6158
rect 6545 6155 6611 6158
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 3233 5946 3299 5949
rect 4153 5946 4219 5949
rect 3233 5944 4219 5946
rect 3233 5888 3238 5944
rect 3294 5888 4158 5944
rect 4214 5888 4219 5944
rect 3233 5886 4219 5888
rect 3233 5883 3299 5886
rect 4153 5883 4219 5886
rect 5809 5946 5875 5949
rect 6729 5946 6795 5949
rect 5809 5944 6795 5946
rect 5809 5888 5814 5944
rect 5870 5888 6734 5944
rect 6790 5888 6795 5944
rect 5809 5886 6795 5888
rect 5809 5883 5875 5886
rect 6729 5883 6795 5886
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 3509 5810 3575 5813
rect 6269 5810 6335 5813
rect 3509 5808 6335 5810
rect 3509 5752 3514 5808
rect 3570 5752 6274 5808
rect 6330 5752 6335 5808
rect 3509 5750 6335 5752
rect 3509 5747 3575 5750
rect 6269 5747 6335 5750
rect 8201 5810 8267 5813
rect 11200 5810 12000 5840
rect 8201 5808 12000 5810
rect 8201 5752 8206 5808
rect 8262 5752 12000 5808
rect 8201 5750 12000 5752
rect 8201 5747 8267 5750
rect 11200 5720 12000 5750
rect 1669 5674 1735 5677
rect 3233 5674 3299 5677
rect 1669 5672 3299 5674
rect 1669 5616 1674 5672
rect 1730 5616 3238 5672
rect 3294 5616 3299 5672
rect 1669 5614 3299 5616
rect 1669 5611 1735 5614
rect 3233 5611 3299 5614
rect 3601 5674 3667 5677
rect 3601 5672 4170 5674
rect 3601 5616 3606 5672
rect 3662 5616 4170 5672
rect 3601 5614 4170 5616
rect 3601 5611 3667 5614
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 3049 5402 3115 5405
rect 3049 5400 3250 5402
rect 3049 5344 3054 5400
rect 3110 5344 3250 5400
rect 3049 5342 3250 5344
rect 3049 5339 3115 5342
rect 1945 5266 2011 5269
rect 1945 5264 3066 5266
rect 1945 5208 1950 5264
rect 2006 5208 3066 5264
rect 1945 5206 3066 5208
rect 1945 5203 2011 5206
rect 2313 5130 2379 5133
rect 2313 5128 2790 5130
rect 2313 5072 2318 5128
rect 2374 5072 2790 5128
rect 2313 5070 2790 5072
rect 2313 5067 2379 5070
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 2730 4586 2790 5070
rect 3006 4994 3066 5206
rect 3190 5130 3250 5342
rect 4110 5266 4170 5614
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 10698 5407 11014 5408
rect 9029 5266 9095 5269
rect 4110 5264 9095 5266
rect 4110 5208 9034 5264
rect 9090 5208 9095 5264
rect 4110 5206 9095 5208
rect 9029 5203 9095 5206
rect 5625 5130 5691 5133
rect 3190 5128 5691 5130
rect 3190 5072 5630 5128
rect 5686 5072 5691 5128
rect 3190 5070 5691 5072
rect 5625 5067 5691 5070
rect 3969 4994 4035 4997
rect 3006 4992 4035 4994
rect 3006 4936 3974 4992
rect 4030 4936 4035 4992
rect 3006 4934 4035 4936
rect 3969 4931 4035 4934
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 6269 4722 6335 4725
rect 9673 4722 9739 4725
rect 11200 4722 12000 4752
rect 6269 4720 9739 4722
rect 6269 4664 6274 4720
rect 6330 4664 9678 4720
rect 9734 4664 9739 4720
rect 6269 4662 9739 4664
rect 6269 4659 6335 4662
rect 9673 4659 9739 4662
rect 10504 4662 12000 4722
rect 2865 4586 2931 4589
rect 2730 4584 2931 4586
rect 2730 4528 2870 4584
rect 2926 4528 2931 4584
rect 2730 4526 2931 4528
rect 2865 4523 2931 4526
rect 3049 4586 3115 4589
rect 10133 4586 10199 4589
rect 3049 4584 10199 4586
rect 3049 4528 3054 4584
rect 3110 4528 10138 4584
rect 10194 4528 10199 4584
rect 3049 4526 10199 4528
rect 3049 4523 3115 4526
rect 10133 4523 10199 4526
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 4337 4314 4403 4317
rect 4797 4314 4863 4317
rect 4337 4312 4863 4314
rect 4337 4256 4342 4312
rect 4398 4256 4802 4312
rect 4858 4256 4863 4312
rect 4337 4254 4863 4256
rect 4337 4251 4403 4254
rect 4797 4251 4863 4254
rect 10504 4178 10564 4662
rect 11200 4632 12000 4662
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 10698 4319 11014 4320
rect 2454 4118 10564 4178
rect 2454 4045 2514 4118
rect 2454 4040 2563 4045
rect 2454 3984 2502 4040
rect 2558 3984 2563 4040
rect 2454 3982 2563 3984
rect 2497 3979 2563 3982
rect 2681 4042 2747 4045
rect 8017 4042 8083 4045
rect 2681 4040 8083 4042
rect 2681 3984 2686 4040
rect 2742 3984 8022 4040
rect 8078 3984 8083 4040
rect 2681 3982 8083 3984
rect 2681 3979 2747 3982
rect 8017 3979 8083 3982
rect 3182 3844 3188 3908
rect 3252 3906 3258 3908
rect 3509 3906 3575 3909
rect 3252 3904 3575 3906
rect 3252 3848 3514 3904
rect 3570 3848 3575 3904
rect 3252 3846 3575 3848
rect 3252 3844 3258 3846
rect 3509 3843 3575 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 0 3634 800 3664
rect 2957 3634 3023 3637
rect 0 3632 3023 3634
rect 0 3576 2962 3632
rect 3018 3576 3023 3632
rect 0 3574 3023 3576
rect 0 3544 800 3574
rect 2957 3571 3023 3574
rect 5073 3634 5139 3637
rect 11200 3634 12000 3664
rect 5073 3632 12000 3634
rect 5073 3576 5078 3632
rect 5134 3576 12000 3632
rect 5073 3574 12000 3576
rect 5073 3571 5139 3574
rect 11200 3544 12000 3574
rect 2405 3498 2471 3501
rect 7281 3498 7347 3501
rect 2405 3496 7347 3498
rect 2405 3440 2410 3496
rect 2466 3440 7286 3496
rect 7342 3440 7347 3496
rect 2405 3438 7347 3440
rect 2405 3435 2471 3438
rect 7281 3435 7347 3438
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 10698 3231 11014 3232
rect 1894 3028 1900 3092
rect 1964 3090 1970 3092
rect 5625 3090 5691 3093
rect 1964 3088 5691 3090
rect 1964 3032 5630 3088
rect 5686 3032 5691 3088
rect 1964 3030 5691 3032
rect 1964 3028 1970 3030
rect 5625 3027 5691 3030
rect 2405 2954 2471 2957
rect 9949 2954 10015 2957
rect 2405 2952 10015 2954
rect 2405 2896 2410 2952
rect 2466 2896 9954 2952
rect 10010 2896 10015 2952
rect 2405 2894 10015 2896
rect 2405 2891 2471 2894
rect 9949 2891 10015 2894
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 0 2546 800 2576
rect 1577 2546 1643 2549
rect 0 2544 1643 2546
rect 0 2488 1582 2544
rect 1638 2488 1643 2544
rect 0 2486 1643 2488
rect 0 2456 800 2486
rect 1577 2483 1643 2486
rect 7465 2546 7531 2549
rect 11200 2546 12000 2576
rect 7465 2544 12000 2546
rect 7465 2488 7470 2544
rect 7526 2488 12000 2544
rect 7465 2486 12000 2488
rect 7465 2483 7531 2486
rect 11200 2456 12000 2486
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 10698 2143 11014 2144
rect 0 1458 800 1488
rect 6729 1458 6795 1461
rect 0 1456 6795 1458
rect 0 1400 6734 1456
rect 6790 1400 6795 1456
rect 0 1398 6795 1400
rect 0 1368 800 1398
rect 6729 1395 6795 1398
rect 8937 1458 9003 1461
rect 11200 1458 12000 1488
rect 8937 1456 12000 1458
rect 8937 1400 8942 1456
rect 8998 1400 12000 1456
rect 8937 1398 12000 1400
rect 8937 1395 9003 1398
rect 11200 1368 12000 1398
rect 9305 370 9371 373
rect 11200 370 12000 400
rect 9305 368 12000 370
rect 9305 312 9310 368
rect 9366 312 12000 368
rect 9305 310 12000 312
rect 9305 307 9371 310
rect 11200 280 12000 310
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 1900 8332 1964 8396
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3188 6700 3252 6764
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 3188 3844 3252 3908
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 1900 3028 1964 3092
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 1899 8396 1965 8397
rect 1899 8332 1900 8396
rect 1964 8332 1965 8396
rect 1899 8331 1965 8332
rect 1902 3093 1962 8331
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3187 6764 3253 6765
rect 3187 6700 3188 6764
rect 3252 6700 3253 6764
rect 3187 6699 3253 6700
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 3190 3909 3250 6699
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3187 3908 3253 3909
rect 3187 3844 3188 3908
rect 3252 3844 3253 3908
rect 3187 3843 3253 3844
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 1899 3092 1965 3093
rect 1899 3028 1900 3092
rect 1964 3028 1965 3092
rect 1899 3027 1965 3028
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform 1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1688980957
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1688980957
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1688980957
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1688980957
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1688980957
transform 1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1688980957
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1688980957
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1688980957
transform 1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1688980957
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1688980957
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 1688980957
transform 1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _119_
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _121_
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _122_
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _123_
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _124_
timestamp 1688980957
transform 1 0 6900 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _125_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _126_
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _127_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1688980957
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _150__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _150_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _151_
timestamp 1688980957
transform 1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _152_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _153_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _154_
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _155_
timestamp 1688980957
transform 1 0 6532 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _156_
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _157_
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _158_
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _159_
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _160_
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _161_
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _162_
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _163_
timestamp 1688980957
transform 1 0 4416 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _163__44
timestamp 1688980957
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _164_
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _165_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _166_
timestamp 1688980957
transform 1 0 2392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _167_
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _168_
timestamp 1688980957
transform 1 0 5428 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _169_
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _170_
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _171_
timestamp 1688980957
transform 1 0 3496 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _172_
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _173_
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _174_
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _174__45
timestamp 1688980957
transform -1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _175_
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _176_
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _177_
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _178__46
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _178_
timestamp 1688980957
transform 1 0 9568 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _179_
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _180_
timestamp 1688980957
transform 1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _181_
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_8
timestamp 1688980957
transform 1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_52
timestamp 1688980957
transform 1 0 5888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_11
timestamp 1688980957
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_56
timestamp 1688980957
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_91
timestamp 1688980957
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_102
timestamp 1688980957
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_12
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_29
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_74
timestamp 1688980957
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_83
timestamp 1688980957
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_40
timestamp 1688980957
transform 1 0 4784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_93
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_11
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_21
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_40
timestamp 1688980957
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_101
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_45
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_91
timestamp 1688980957
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_101
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_28
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_46
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_101
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_8
timestamp 1688980957
transform 1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_59
timestamp 1688980957
transform 1 0 6532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_98
timestamp 1688980957
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_50
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_56
timestamp 1688980957
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_74
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_82
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_40
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_57
timestamp 1688980957
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1688980957
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_6
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_20
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_40
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_46
timestamp 1688980957
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_66
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_72
timestamp 1688980957
transform 1 0 7728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1688980957
transform 1 0 1840 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform 1 0 5428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform 1 0 6624 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 6532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
port 0 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
port 1 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
port 2 nsew signal tristate
flabel metal3 s 11200 10072 12000 10192 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 11200 11160 12000 11280 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 5 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 6 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 7 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 8 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 9 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 10 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 11 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 12 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 13 nsew signal input
flabel metal2 s 570 11200 626 12000 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 14 nsew signal tristate
flabel metal2 s 1766 11200 1822 12000 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 15 nsew signal tristate
flabel metal2 s 2962 11200 3018 12000 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 16 nsew signal tristate
flabel metal2 s 4158 11200 4214 12000 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 17 nsew signal tristate
flabel metal2 s 5354 11200 5410 12000 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 18 nsew signal tristate
flabel metal2 s 6550 11200 6606 12000 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 19 nsew signal tristate
flabel metal2 s 7746 11200 7802 12000 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 20 nsew signal tristate
flabel metal2 s 8942 11200 8998 12000 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 21 nsew signal tristate
flabel metal2 s 10138 11200 10194 12000 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 22 nsew signal tristate
flabel metal3 s 11200 280 12000 400 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 23 nsew signal input
flabel metal3 s 11200 1368 12000 1488 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 24 nsew signal input
flabel metal3 s 11200 2456 12000 2576 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 25 nsew signal input
flabel metal3 s 11200 3544 12000 3664 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 26 nsew signal input
flabel metal3 s 11200 4632 12000 4752 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 27 nsew signal input
flabel metal3 s 11200 5720 12000 5840 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 28 nsew signal input
flabel metal3 s 11200 6808 12000 6928 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 29 nsew signal input
flabel metal3 s 11200 7896 12000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 30 nsew signal input
flabel metal3 s 11200 8984 12000 9104 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 31 nsew signal input
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 32 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 33 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 34 nsew signal tristate
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 35 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 36 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 37 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 38 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 39 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 40 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 41 nsew signal input
flabel metal2 s 11334 11200 11390 12000 0 FreeSans 224 90 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
port 42 nsew signal tristate
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 4370 3366 4370 3366 0 _000_
rlabel metal1 3450 5712 3450 5712 0 _001_
rlabel metal2 2898 6426 2898 6426 0 _002_
rlabel metal1 6302 6426 6302 6426 0 _003_
rlabel metal1 5106 7412 5106 7412 0 _004_
rlabel metal1 9522 6256 9522 6256 0 _005_
rlabel metal1 9706 7514 9706 7514 0 _006_
rlabel metal1 5566 5202 5566 5202 0 _007_
rlabel metal1 8832 6290 8832 6290 0 _008_
rlabel metal1 9660 5882 9660 5882 0 _009_
rlabel metal1 6578 5678 6578 5678 0 _010_
rlabel metal1 7222 2482 7222 2482 0 _011_
rlabel metal1 8740 3366 8740 3366 0 _012_
rlabel metal1 4600 5066 4600 5066 0 _013_
rlabel metal2 2806 6324 2806 6324 0 _014_
rlabel metal1 2300 4114 2300 4114 0 _015_
rlabel metal1 8280 6426 8280 6426 0 _016_
rlabel metal1 6348 4658 6348 4658 0 _017_
rlabel metal2 9338 6936 9338 6936 0 _018_
rlabel metal1 5658 7276 5658 7276 0 _019_
rlabel metal1 10074 7922 10074 7922 0 _020_
rlabel metal1 6578 7378 6578 7378 0 _021_
rlabel metal1 5750 5100 5750 5100 0 _022_
rlabel metal1 6164 5882 6164 5882 0 _023_
rlabel metal1 7452 6970 7452 6970 0 _024_
rlabel metal1 7130 5746 7130 5746 0 _025_
rlabel metal1 7452 7922 7452 7922 0 _026_
rlabel metal2 9706 6528 9706 6528 0 _027_
rlabel metal1 6118 2278 6118 2278 0 _028_
rlabel metal2 4646 3604 4646 3604 0 _029_
rlabel metal2 2622 5389 2622 5389 0 _030_
rlabel metal1 3956 5678 3956 5678 0 _031_
rlabel metal2 1978 4454 1978 4454 0 _032_
rlabel metal1 5796 4590 5796 4590 0 _033_
rlabel metal2 3082 5899 3082 5899 0 _034_
rlabel metal1 4584 4114 4584 4114 0 _035_
rlabel metal2 1978 5933 1978 5933 0 _036_
rlabel metal1 4186 4794 4186 4794 0 _037_
rlabel metal1 2346 2516 2346 2516 0 _038_
rlabel metal1 4232 4046 4232 4046 0 _039_
rlabel metal2 9890 3723 9890 3723 0 _040_
rlabel metal1 7314 2550 7314 2550 0 _041_
rlabel metal2 9154 2210 9154 2210 0 _042_
rlabel metal1 8004 2482 8004 2482 0 _043_
rlabel metal2 8280 5610 8280 5610 0 _044_
rlabel metal2 9890 5100 9890 5100 0 _045_
rlabel metal1 9982 4488 9982 4488 0 _046_
rlabel metal1 8096 5678 8096 5678 0 _047_
rlabel metal2 8694 1639 8694 1639 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_
rlabel metal2 9614 1520 9614 1520 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_
rlabel metal1 10442 2958 10442 2958 0 bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_
rlabel metal1 8786 9622 8786 9622 0 ccff_head
rlabel metal1 9798 9146 9798 9146 0 ccff_tail
rlabel metal3 1142 2516 1142 2516 0 chanx_left_in[0]
rlabel metal3 1832 3604 1832 3604 0 chanx_left_in[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_in[2]
rlabel metal3 820 5780 820 5780 0 chanx_left_in[3]
rlabel metal3 1050 6868 1050 6868 0 chanx_left_in[4]
rlabel metal3 751 7956 751 7956 0 chanx_left_in[5]
rlabel metal3 820 9044 820 9044 0 chanx_left_in[6]
rlabel metal3 1740 10132 1740 10132 0 chanx_left_in[7]
rlabel metal3 1027 11220 1027 11220 0 chanx_left_in[8]
rlabel metal1 1104 9146 1104 9146 0 chanx_left_out[0]
rlabel metal1 2070 9622 2070 9622 0 chanx_left_out[1]
rlabel metal1 3266 9622 3266 9622 0 chanx_left_out[2]
rlabel metal1 4462 9622 4462 9622 0 chanx_left_out[3]
rlabel metal1 5566 9418 5566 9418 0 chanx_left_out[4]
rlabel metal1 6716 9690 6716 9690 0 chanx_left_out[5]
rlabel metal1 7958 9418 7958 9418 0 chanx_left_out[6]
rlabel metal1 9246 9622 9246 9622 0 chanx_left_out[7]
rlabel metal1 10258 9418 10258 9418 0 chanx_left_out[8]
rlabel metal1 10350 2448 10350 2448 0 chanx_right_in[0]
rlabel metal2 8924 1428 8924 1428 0 chanx_right_in[1]
rlabel metal3 9392 2516 9392 2516 0 chanx_right_in[2]
rlabel metal1 3910 3468 3910 3468 0 chanx_right_in[3]
rlabel metal1 2070 3060 2070 3060 0 chanx_right_in[4]
rlabel metal1 9154 7854 9154 7854 0 chanx_right_in[5]
rlabel metal1 10718 7378 10718 7378 0 chanx_right_in[6]
rlabel metal1 9798 8432 9798 8432 0 chanx_right_in[7]
rlabel metal1 9798 9588 9798 9588 0 chanx_right_in[8]
rlabel metal1 1012 3910 1012 3910 0 chanx_right_out[0]
rlabel metal1 1472 4454 1472 4454 0 chanx_right_out[1]
rlabel metal2 2254 959 2254 959 0 chanx_right_out[2]
rlabel metal2 3174 1520 3174 1520 0 chanx_right_out[3]
rlabel metal2 4094 959 4094 959 0 chanx_right_out[4]
rlabel metal2 5014 1520 5014 1520 0 chanx_right_out[5]
rlabel metal2 5934 823 5934 823 0 chanx_right_out[6]
rlabel metal2 6854 1095 6854 1095 0 chanx_right_out[7]
rlabel metal2 7774 1095 7774 1095 0 chanx_right_out[8]
rlabel metal1 2691 3094 2691 3094 0 clknet_0_prog_clk
rlabel metal1 2346 3978 2346 3978 0 clknet_1_0__leaf_prog_clk
rlabel metal1 8418 5236 8418 5236 0 clknet_1_1__leaf_prog_clk
rlabel metal1 10350 6664 10350 6664 0 mem_bottom_ipin_0.DFF_0_.Q
rlabel metal1 6762 7854 6762 7854 0 mem_bottom_ipin_0.DFF_1_.Q
rlabel metal1 7912 6086 7912 6086 0 mem_bottom_ipin_0.DFF_2_.Q
rlabel metal1 2530 6732 2530 6732 0 mem_top_ipin_0.DFF_0_.Q
rlabel metal1 1978 6766 1978 6766 0 mem_top_ipin_0.DFF_1_.Q
rlabel metal1 5842 4046 5842 4046 0 mem_top_ipin_0.DFF_2_.Q
rlabel metal1 6946 4114 6946 4114 0 mem_top_ipin_1.DFF_0_.Q
rlabel metal2 2714 3757 2714 3757 0 mem_top_ipin_1.DFF_1_.Q
rlabel metal1 9430 5712 9430 5712 0 mem_top_ipin_2.DFF_0_.Q
rlabel metal1 4048 4658 4048 4658 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 6532 4590 6532 4590 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 4278 6766 4278 6766 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal1 5382 7310 5382 7310 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 7130 7854 7130 7854 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal1 9522 7922 9522 7922 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal2 6946 5202 6946 5202 0 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 5842 6970 5842 6970 0 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 8924 7990 8924 7990 0 mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 7820 6834 7820 6834 0 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8418 7480 8418 7480 0 mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 9154 7310 9154 7310 0 mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 2070 2482 2070 2482 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 2438 4556 2438 4556 0 mux_top_ipin_0.INVTX1_3_.out
rlabel metal1 3450 5134 3450 5134 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal1 4232 5338 4232 5338 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal1 5796 4726 5796 4726 0 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2852 3570 2852 3570 0 mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4462 5270 4462 5270 0 mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 5566 3400 5566 3400 0 mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 5014 3808 5014 3808 0 mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 6164 3638 6164 3638 0 mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 7728 2482 7728 2482 0 mux_top_ipin_1.INVTX1_0_.out
rlabel metal1 4945 2550 4945 2550 0 mux_top_ipin_1.INVTX1_1_.out
rlabel metal1 8004 2550 8004 2550 0 mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9936 2550 9936 2550 0 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8556 5746 8556 5746 0 mux_top_ipin_2.INVTX1_0_.out
rlabel via2 2438 2907 2438 2907 0 mux_top_ipin_2.INVTX1_1_.out
rlabel metal1 9890 4692 9890 4692 0 mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 10166 4692 10166 4692 0 mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9144 6766 9144 6766 0 net1
rlabel metal1 6946 7820 6946 7820 0 net10
rlabel metal1 7130 2312 7130 2312 0 net11
rlabel metal1 2162 8942 2162 8942 0 net12
rlabel metal2 2346 5389 2346 5389 0 net13
rlabel metal1 4140 3706 4140 3706 0 net14
rlabel metal1 1840 3162 1840 3162 0 net15
rlabel metal1 5658 6324 5658 6324 0 net16
rlabel metal1 10212 7378 10212 7378 0 net17
rlabel metal1 9568 8466 9568 8466 0 net18
rlabel metal1 9706 8942 9706 8942 0 net19
rlabel metal1 2300 4590 2300 4590 0 net2
rlabel metal1 9706 5202 9706 5202 0 net20
rlabel metal2 10028 2346 10028 2346 0 net21
rlabel metal1 6486 3536 6486 3536 0 net22
rlabel metal2 9246 8636 9246 8636 0 net23
rlabel metal4 1932 5712 1932 5712 0 net24
rlabel metal1 2024 9146 2024 9146 0 net25
rlabel metal1 2438 5542 2438 5542 0 net26
rlabel metal1 4462 9146 4462 9146 0 net27
rlabel metal1 5520 8058 5520 8058 0 net28
rlabel metal1 5612 6426 5612 6426 0 net29
rlabel metal1 1610 5644 1610 5644 0 net3
rlabel metal1 9982 7242 9982 7242 0 net30
rlabel metal1 9246 8602 9246 8602 0 net31
rlabel metal2 9246 9316 9246 9316 0 net32
rlabel metal1 1840 4182 1840 4182 0 net33
rlabel metal1 1518 4658 1518 4658 0 net34
rlabel metal1 1702 2380 1702 2380 0 net35
rlabel metal2 3266 4029 3266 4029 0 net36
rlabel metal1 3818 2414 3818 2414 0 net37
rlabel metal1 5106 2414 5106 2414 0 net38
rlabel metal1 7360 4182 7360 4182 0 net39
rlabel metal1 2254 5236 2254 5236 0 net4
rlabel metal1 6394 8806 6394 8806 0 net40
rlabel metal1 10028 3094 10028 3094 0 net41
rlabel metal1 9936 8602 9936 8602 0 net42
rlabel metal1 7636 7378 7636 7378 0 net43
rlabel metal1 4186 2482 4186 2482 0 net44
rlabel via2 2438 3451 2438 3451 0 net45
rlabel metal1 9706 5780 9706 5780 0 net46
rlabel metal1 6849 3026 6849 3026 0 net47
rlabel metal1 6762 5882 6762 5882 0 net48
rlabel metal1 9154 4794 9154 4794 0 net49
rlabel metal1 1886 6324 1886 6324 0 net5
rlabel metal1 7585 3502 7585 3502 0 net50
rlabel metal2 8694 4386 8694 4386 0 net51
rlabel metal1 7079 6290 7079 6290 0 net52
rlabel metal1 8096 6154 8096 6154 0 net53
rlabel metal1 3910 4148 3910 4148 0 net54
rlabel metal1 4630 3094 4630 3094 0 net55
rlabel metal1 2484 6290 2484 6290 0 net6
rlabel metal1 2254 6256 2254 6256 0 net7
rlabel metal1 1426 8568 1426 8568 0 net8
rlabel metal2 2714 9248 2714 9248 0 net9
rlabel metal3 3718 1428 3718 1428 0 prog_clk
rlabel metal1 10028 8874 10028 8874 0 top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
