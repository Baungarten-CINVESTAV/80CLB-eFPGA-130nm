magic
tech sky130A
magscale 1 2
timestamp 1708041460
<< viali >>
rect 13829 17289 13863 17323
rect 2789 17221 2823 17255
rect 1869 17153 1903 17187
rect 2421 17153 2455 17187
rect 13553 17153 13587 17187
rect 14473 17153 14507 17187
rect 1961 16949 1995 16983
rect 14289 16949 14323 16983
rect 1777 16745 1811 16779
rect 2237 16745 2271 16779
rect 2145 16541 2179 16575
rect 8401 16541 8435 16575
rect 13921 16541 13955 16575
rect 14289 16541 14323 16575
rect 1685 16473 1719 16507
rect 8217 16405 8251 16439
rect 13737 16405 13771 16439
rect 14473 16405 14507 16439
rect 1593 16201 1627 16235
rect 1501 16065 1535 16099
rect 2145 15657 2179 15691
rect 14381 15657 14415 15691
rect 1501 15453 1535 15487
rect 5641 15453 5675 15487
rect 14197 15453 14231 15487
rect 2053 15385 2087 15419
rect 1593 15317 1627 15351
rect 5733 15317 5767 15351
rect 2605 15045 2639 15079
rect 1593 14977 1627 15011
rect 2237 14977 2271 15011
rect 2513 14977 2547 15011
rect 2789 14977 2823 15011
rect 2881 14977 2915 15011
rect 3065 14977 3099 15011
rect 14197 14977 14231 15011
rect 2421 14841 2455 14875
rect 1409 14773 1443 14807
rect 1961 14773 1995 14807
rect 3249 14773 3283 14807
rect 14381 14773 14415 14807
rect 1777 14501 1811 14535
rect 10057 14501 10091 14535
rect 2421 14433 2455 14467
rect 1961 14365 1995 14399
rect 2237 14365 2271 14399
rect 2329 14365 2363 14399
rect 2881 14365 2915 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 8585 14365 8619 14399
rect 10425 14365 10459 14399
rect 10701 14365 10735 14399
rect 9505 14297 9539 14331
rect 9597 14297 9631 14331
rect 1685 14229 1719 14263
rect 2053 14229 2087 14263
rect 3341 14229 3375 14263
rect 3617 14229 3651 14263
rect 4077 14229 4111 14263
rect 8401 14229 8435 14263
rect 8953 14229 8987 14263
rect 10241 14229 10275 14263
rect 10517 14229 10551 14263
rect 2881 14025 2915 14059
rect 3433 14025 3467 14059
rect 3893 14025 3927 14059
rect 8585 14025 8619 14059
rect 1501 13957 1535 13991
rect 2789 13957 2823 13991
rect 9689 13957 9723 13991
rect 10425 13957 10459 13991
rect 1961 13889 1995 13923
rect 2237 13889 2271 13923
rect 2329 13889 2363 13923
rect 3065 13889 3099 13923
rect 3341 13889 3375 13923
rect 3617 13889 3651 13923
rect 3709 13889 3743 13923
rect 3985 13889 4019 13923
rect 4077 13889 4111 13923
rect 4445 13889 4479 13923
rect 4721 13889 4755 13923
rect 10333 13889 10367 13923
rect 12633 13889 12667 13923
rect 14105 13889 14139 13923
rect 2053 13821 2087 13855
rect 7941 13821 7975 13855
rect 8125 13821 8159 13855
rect 8677 13821 8711 13855
rect 9597 13821 9631 13855
rect 9873 13821 9907 13855
rect 14381 13821 14415 13855
rect 4261 13753 4295 13787
rect 1593 13685 1627 13719
rect 3157 13685 3191 13719
rect 9321 13685 9355 13719
rect 12725 13685 12759 13719
rect 3065 13481 3099 13515
rect 7757 13481 7791 13515
rect 8585 13481 8619 13515
rect 10333 13481 10367 13515
rect 13921 13481 13955 13515
rect 7389 13413 7423 13447
rect 2513 13345 2547 13379
rect 8125 13345 8159 13379
rect 12817 13345 12851 13379
rect 2145 13277 2179 13311
rect 2421 13277 2455 13311
rect 2881 13277 2915 13311
rect 3157 13277 3191 13311
rect 3433 13277 3467 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 5089 13277 5123 13311
rect 7573 13277 7607 13311
rect 7665 13277 7699 13311
rect 7941 13277 7975 13311
rect 8953 13277 8987 13311
rect 11253 13277 11287 13311
rect 11520 13277 11554 13311
rect 13001 13277 13035 13311
rect 13737 13277 13771 13311
rect 14197 13277 14231 13311
rect 1501 13209 1535 13243
rect 9220 13209 9254 13243
rect 1593 13141 1627 13175
rect 2329 13141 2363 13175
rect 3341 13141 3375 13175
rect 3617 13141 3651 13175
rect 4997 13141 5031 13175
rect 5181 13141 5215 13175
rect 12633 13141 12667 13175
rect 13461 13141 13495 13175
rect 14381 13141 14415 13175
rect 3525 12937 3559 12971
rect 8309 12937 8343 12971
rect 12357 12937 12391 12971
rect 13553 12937 13587 12971
rect 3985 12869 4019 12903
rect 4997 12869 5031 12903
rect 5549 12869 5583 12903
rect 1777 12801 1811 12835
rect 1869 12801 1903 12835
rect 2881 12801 2915 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 7012 12801 7046 12835
rect 8493 12801 8527 12835
rect 9229 12801 9263 12835
rect 9505 12801 9539 12835
rect 10333 12801 10367 12835
rect 11069 12801 11103 12835
rect 11345 12801 11379 12835
rect 12265 12801 12299 12835
rect 13001 12801 13035 12835
rect 13277 12801 13311 12835
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 14105 12801 14139 12835
rect 2329 12733 2363 12767
rect 3065 12733 3099 12767
rect 3893 12733 3927 12767
rect 4169 12733 4203 12767
rect 5825 12733 5859 12767
rect 6745 12733 6779 12767
rect 8585 12733 8619 12767
rect 8769 12733 8803 12767
rect 1961 12665 1995 12699
rect 8125 12665 8159 12699
rect 9321 12665 9355 12699
rect 10885 12665 10919 12699
rect 13829 12665 13863 12699
rect 1593 12597 1627 12631
rect 2697 12597 2731 12631
rect 5181 12597 5215 12631
rect 10149 12597 10183 12631
rect 11161 12597 11195 12631
rect 13185 12597 13219 12631
rect 13461 12597 13495 12631
rect 14197 12597 14231 12631
rect 2605 12393 2639 12427
rect 7297 12393 7331 12427
rect 7389 12393 7423 12427
rect 9321 12393 9355 12427
rect 12909 12393 12943 12427
rect 13737 12393 13771 12427
rect 6285 12325 6319 12359
rect 10701 12325 10735 12359
rect 11161 12325 11195 12359
rect 14381 12325 14415 12359
rect 4445 12257 4479 12291
rect 7665 12257 7699 12291
rect 7849 12257 7883 12291
rect 9137 12257 9171 12291
rect 9781 12257 9815 12291
rect 10793 12257 10827 12291
rect 11529 12257 11563 12291
rect 12173 12257 12207 12291
rect 12449 12257 12483 12291
rect 13001 12257 13035 12291
rect 2145 12189 2179 12223
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 3985 12189 4019 12223
rect 4905 12189 4939 12223
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 7573 12189 7607 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9689 12189 9723 12223
rect 10057 12189 10091 12223
rect 10241 12189 10275 12223
rect 10977 12189 11011 12223
rect 12265 12189 12299 12223
rect 13185 12189 13219 12223
rect 13921 12189 13955 12223
rect 14197 12189 14231 12223
rect 1501 12121 1535 12155
rect 4169 12121 4203 12155
rect 4261 12121 4295 12155
rect 5172 12121 5206 12155
rect 1593 12053 1627 12087
rect 1961 12053 1995 12087
rect 3617 12053 3651 12087
rect 3801 12053 3835 12087
rect 6469 12053 6503 12087
rect 8309 12053 8343 12087
rect 8493 12053 8527 12087
rect 13645 12053 13679 12087
rect 2145 11849 2179 11883
rect 2605 11849 2639 11883
rect 4445 11849 4479 11883
rect 5365 11849 5399 11883
rect 7113 11849 7147 11883
rect 8309 11849 8343 11883
rect 9965 11849 9999 11883
rect 10333 11849 10367 11883
rect 11989 11849 12023 11883
rect 12265 11849 12299 11883
rect 13645 11849 13679 11883
rect 14013 11849 14047 11883
rect 1869 11781 1903 11815
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 2053 11713 2087 11747
rect 2329 11713 2363 11747
rect 2789 11713 2823 11747
rect 3148 11713 3182 11747
rect 4629 11713 4663 11747
rect 4721 11713 4755 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 7573 11713 7607 11747
rect 7849 11713 7883 11747
rect 10149 11713 10183 11747
rect 10241 11713 10275 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 12541 11713 12575 11747
rect 12633 11713 12667 11747
rect 13185 11713 13219 11747
rect 13921 11713 13955 11747
rect 14197 11713 14231 11747
rect 2881 11645 2915 11679
rect 5457 11645 5491 11679
rect 6561 11645 6595 11679
rect 7665 11645 7699 11679
rect 13001 11645 13035 11679
rect 4261 11577 4295 11611
rect 6837 11577 6871 11611
rect 1501 11509 1535 11543
rect 2421 11509 2455 11543
rect 6101 11509 6135 11543
rect 7389 11509 7423 11543
rect 11713 11509 11747 11543
rect 14381 11509 14415 11543
rect 1409 11305 1443 11339
rect 2973 11305 3007 11339
rect 3433 11305 3467 11339
rect 9321 11305 9355 11339
rect 11897 11305 11931 11339
rect 1869 11237 1903 11271
rect 4169 11237 4203 11271
rect 7665 11237 7699 11271
rect 7849 11237 7883 11271
rect 8125 11237 8159 11271
rect 14105 11237 14139 11271
rect 2421 11169 2455 11203
rect 3249 11169 3283 11203
rect 3985 11169 4019 11203
rect 6285 11169 6319 11203
rect 9137 11169 9171 11203
rect 11989 11169 12023 11203
rect 13093 11169 13127 11203
rect 1593 11101 1627 11135
rect 1685 11101 1719 11135
rect 1961 11101 1995 11135
rect 3157 11101 3191 11135
rect 3617 11101 3651 11135
rect 3801 11101 3835 11135
rect 4721 11101 4755 11135
rect 6469 11101 6503 11135
rect 8033 11101 8067 11135
rect 8309 11101 8343 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 10517 11101 10551 11135
rect 12725 11101 12759 11135
rect 14289 11101 14323 11135
rect 4988 11033 5022 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 7205 11033 7239 11067
rect 10784 11033 10818 11067
rect 13185 11033 13219 11067
rect 13737 11033 13771 11067
rect 6101 10965 6135 10999
rect 8493 10965 8527 10999
rect 12633 10965 12667 10999
rect 12817 10965 12851 10999
rect 2881 10761 2915 10795
rect 5181 10761 5215 10795
rect 5273 10761 5307 10795
rect 7849 10761 7883 10795
rect 8493 10761 8527 10795
rect 9321 10761 9355 10795
rect 13461 10761 13495 10795
rect 6193 10693 6227 10727
rect 6561 10693 6595 10727
rect 11888 10693 11922 10727
rect 13921 10693 13955 10727
rect 1593 10625 1627 10659
rect 1961 10625 1995 10659
rect 3065 10625 3099 10659
rect 3157 10625 3191 10659
rect 3617 10625 3651 10659
rect 3801 10625 3835 10659
rect 4068 10625 4102 10659
rect 5457 10625 5491 10659
rect 7113 10625 7147 10659
rect 7941 10625 7975 10659
rect 8401 10625 8435 10659
rect 8861 10625 8895 10659
rect 9413 10625 9447 10659
rect 10149 10625 10183 10659
rect 10609 10625 10643 10659
rect 11621 10625 11655 10659
rect 13645 10625 13679 10659
rect 2145 10557 2179 10591
rect 2329 10557 2363 10591
rect 5641 10557 5675 10591
rect 6469 10557 6503 10591
rect 7205 10557 7239 10591
rect 7389 10557 7423 10591
rect 8677 10557 8711 10591
rect 9597 10557 9631 10591
rect 10241 10557 10275 10591
rect 10701 10557 10735 10591
rect 10885 10557 10919 10591
rect 13829 10557 13863 10591
rect 14105 10557 14139 10591
rect 1777 10489 1811 10523
rect 2789 10489 2823 10523
rect 8125 10489 8159 10523
rect 1409 10421 1443 10455
rect 3249 10421 3283 10455
rect 3433 10421 3467 10455
rect 10057 10421 10091 10455
rect 10425 10421 10459 10455
rect 11345 10421 11379 10455
rect 13001 10421 13035 10455
rect 4169 10217 4203 10251
rect 5181 10217 5215 10251
rect 6837 10217 6871 10251
rect 10149 10217 10183 10251
rect 10517 10217 10551 10251
rect 11897 10217 11931 10251
rect 14381 10217 14415 10251
rect 7113 10149 7147 10183
rect 9505 10149 9539 10183
rect 11437 10149 11471 10183
rect 12909 10149 12943 10183
rect 13461 10149 13495 10183
rect 1501 10081 1535 10115
rect 3157 10081 3191 10115
rect 3985 10081 4019 10115
rect 4721 10081 4755 10115
rect 6009 10081 6043 10115
rect 9229 10081 9263 10115
rect 9781 10081 9815 10115
rect 11529 10081 11563 10115
rect 12265 10081 12299 10115
rect 12449 10081 12483 10115
rect 13277 10081 13311 10115
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3801 10013 3835 10047
rect 4537 10013 4571 10047
rect 5365 10013 5399 10047
rect 6193 10013 6227 10047
rect 6745 10013 6779 10047
rect 7021 10013 7055 10047
rect 7297 10013 7331 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 9965 10013 9999 10047
rect 10701 10013 10735 10047
rect 10885 10013 10919 10047
rect 11713 10013 11747 10047
rect 13093 10013 13127 10047
rect 14197 10013 14231 10047
rect 1768 9945 1802 9979
rect 7564 9945 7598 9979
rect 2881 9877 2915 9911
rect 3433 9877 3467 9911
rect 5917 9877 5951 9911
rect 6653 9877 6687 9911
rect 8677 9877 8711 9911
rect 1593 9673 1627 9707
rect 1777 9673 1811 9707
rect 4629 9673 4663 9707
rect 6009 9673 6043 9707
rect 7481 9673 7515 9707
rect 9781 9673 9815 9707
rect 11713 9673 11747 9707
rect 12173 9673 12207 9707
rect 13001 9673 13035 9707
rect 14197 9673 14231 9707
rect 5917 9605 5951 9639
rect 7297 9605 7331 9639
rect 13369 9605 13403 9639
rect 1501 9537 1535 9571
rect 1961 9537 1995 9571
rect 2421 9537 2455 9571
rect 3617 9537 3651 9571
rect 3893 9537 3927 9571
rect 3985 9537 4019 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5457 9537 5491 9571
rect 6201 9537 6235 9571
rect 6561 9537 6595 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 7665 9537 7699 9571
rect 7757 9537 7791 9571
rect 8493 9537 8527 9571
rect 8861 9537 8895 9571
rect 9681 9537 9715 9571
rect 9965 9537 9999 9571
rect 10057 9537 10091 9571
rect 10149 9537 10183 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11161 9537 11195 9571
rect 11621 9537 11655 9571
rect 11897 9537 11931 9571
rect 12357 9537 12391 9571
rect 12633 9537 12667 9571
rect 12909 9537 12943 9571
rect 13277 9537 13311 9571
rect 13737 9537 13771 9571
rect 14105 9537 14139 9571
rect 14381 9537 14415 9571
rect 2513 9469 2547 9503
rect 2697 9469 2731 9503
rect 4169 9469 4203 9503
rect 5273 9469 5307 9503
rect 8217 9469 8251 9503
rect 10333 9469 10367 9503
rect 2237 9401 2271 9435
rect 3433 9401 3467 9435
rect 3709 9401 3743 9435
rect 4721 9401 4755 9435
rect 6377 9401 6411 9435
rect 7113 9401 7147 9435
rect 8585 9401 8619 9435
rect 9505 9401 9539 9435
rect 10609 9401 10643 9435
rect 12449 9401 12483 9435
rect 3157 9333 3191 9367
rect 6745 9333 6779 9367
rect 7941 9333 7975 9367
rect 9413 9333 9447 9367
rect 10977 9333 11011 9367
rect 11253 9333 11287 9367
rect 11989 9333 12023 9367
rect 12725 9333 12759 9367
rect 2145 9129 2179 9163
rect 3065 9129 3099 9163
rect 4261 9129 4295 9163
rect 4997 9129 5031 9163
rect 5733 9129 5767 9163
rect 7205 9129 7239 9163
rect 5273 9061 5307 9095
rect 6101 9061 6135 9095
rect 10333 9061 10367 9095
rect 14381 9061 14415 9095
rect 3525 8993 3559 9027
rect 3985 8993 4019 9027
rect 6469 8993 6503 9027
rect 6653 8993 6687 9027
rect 6837 8993 6871 9027
rect 10517 8993 10551 9027
rect 11989 8993 12023 9027
rect 12173 8993 12207 9027
rect 1593 8925 1627 8959
rect 1869 8925 1903 8959
rect 2329 8925 2363 8959
rect 2605 8925 2639 8959
rect 2697 8925 2731 8959
rect 2882 8925 2916 8959
rect 3433 8925 3467 8959
rect 3801 8925 3835 8959
rect 4721 8925 4755 8959
rect 4813 8925 4847 8959
rect 5089 8925 5123 8959
rect 5365 8925 5399 8959
rect 5641 8925 5675 8959
rect 6285 8925 6319 8959
rect 6377 8925 6411 8959
rect 7389 8925 7423 8959
rect 8953 8925 8987 8959
rect 11253 8925 11287 8959
rect 12817 8925 12851 8959
rect 13645 8925 13679 8959
rect 13737 8925 13771 8959
rect 14197 8925 14231 8959
rect 7656 8857 7690 8891
rect 9220 8857 9254 8891
rect 10609 8857 10643 8891
rect 11161 8857 11195 8891
rect 1409 8789 1443 8823
rect 2053 8789 2087 8823
rect 2421 8789 2455 8823
rect 4537 8789 4571 8823
rect 5457 8789 5491 8823
rect 8769 8789 8803 8823
rect 11897 8789 11931 8823
rect 12633 8789 12667 8823
rect 13369 8789 13403 8823
rect 13461 8789 13495 8823
rect 13921 8789 13955 8823
rect 3433 8585 3467 8619
rect 4169 8585 4203 8619
rect 6377 8585 6411 8619
rect 7297 8585 7331 8619
rect 9689 8585 9723 8619
rect 10885 8585 10919 8619
rect 12909 8585 12943 8619
rect 14473 8585 14507 8619
rect 4804 8517 4838 8551
rect 7389 8517 7423 8551
rect 10057 8517 10091 8551
rect 10149 8517 10183 8551
rect 11796 8517 11830 8551
rect 13093 8517 13127 8551
rect 13185 8517 13219 8551
rect 1777 8449 1811 8483
rect 2605 8449 2639 8483
rect 3525 8449 3559 8483
rect 4261 8449 4295 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 9413 8449 9447 8483
rect 9873 8449 9907 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 11529 8449 11563 8483
rect 13829 8449 13863 8483
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 2881 8381 2915 8415
rect 3709 8381 3743 8415
rect 4537 8381 4571 8415
rect 6653 8381 6687 8415
rect 14013 8381 14047 8415
rect 1593 8313 1627 8347
rect 10609 8313 10643 8347
rect 13645 8313 13679 8347
rect 4353 8245 4387 8279
rect 5917 8245 5951 8279
rect 8677 8245 8711 8279
rect 9229 8245 9263 8279
rect 11345 8245 11379 8279
rect 2237 8041 2271 8075
rect 2697 8041 2731 8075
rect 3617 8041 3651 8075
rect 5181 8041 5215 8075
rect 9229 8041 9263 8075
rect 14197 8041 14231 8075
rect 2421 7973 2455 8007
rect 3157 7905 3191 7939
rect 4445 7905 4479 7939
rect 4997 7905 5031 7939
rect 6837 7905 6871 7939
rect 7021 7905 7055 7939
rect 9413 7905 9447 7939
rect 13093 7905 13127 7939
rect 1409 7837 1443 7871
rect 1869 7837 1903 7871
rect 2145 7837 2179 7871
rect 2605 7837 2639 7871
rect 2881 7837 2915 7871
rect 2973 7837 3007 7871
rect 3801 7837 3835 7871
rect 5089 7837 5123 7871
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 7665 7837 7699 7871
rect 8309 7837 8343 7871
rect 9045 7837 9079 7871
rect 10057 7837 10091 7871
rect 11529 7837 11563 7871
rect 11796 7837 11830 7871
rect 14105 7837 14139 7871
rect 1501 7769 1535 7803
rect 6009 7769 6043 7803
rect 6745 7769 6779 7803
rect 7481 7769 7515 7803
rect 8585 7769 8619 7803
rect 9965 7769 9999 7803
rect 10302 7769 10336 7803
rect 13185 7769 13219 7803
rect 13737 7769 13771 7803
rect 1685 7701 1719 7735
rect 3893 7701 3927 7735
rect 4077 7701 4111 7735
rect 8217 7701 8251 7735
rect 8401 7701 8435 7735
rect 11437 7701 11471 7735
rect 12909 7701 12943 7735
rect 1961 7497 1995 7531
rect 9321 7497 9355 7531
rect 6561 7429 6595 7463
rect 7297 7429 7331 7463
rect 7849 7429 7883 7463
rect 11713 7429 11747 7463
rect 1777 7361 1811 7395
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 2605 7361 2639 7395
rect 4629 7361 4663 7395
rect 5181 7361 5215 7395
rect 6009 7361 6043 7395
rect 7205 7361 7239 7395
rect 7665 7361 7699 7395
rect 9956 7361 9990 7395
rect 11345 7361 11379 7395
rect 13553 7361 13587 7395
rect 14289 7361 14323 7395
rect 4445 7293 4479 7327
rect 5365 7293 5399 7327
rect 6469 7293 6503 7327
rect 9689 7293 9723 7327
rect 11621 7293 11655 7327
rect 12357 7293 12391 7327
rect 12725 7293 12759 7327
rect 13369 7293 13403 7327
rect 1593 7225 1627 7259
rect 3893 7225 3927 7259
rect 5089 7225 5123 7259
rect 5549 7225 5583 7259
rect 7021 7225 7055 7259
rect 7481 7225 7515 7259
rect 12173 7225 12207 7259
rect 2421 7157 2455 7191
rect 6101 7157 6135 7191
rect 11069 7157 11103 7191
rect 11161 7157 11195 7191
rect 13277 7157 13311 7191
rect 13921 7157 13955 7191
rect 14105 7157 14139 7191
rect 3525 6953 3559 6987
rect 5457 6953 5491 6987
rect 13461 6953 13495 6987
rect 6377 6885 6411 6919
rect 5825 6817 5859 6851
rect 6561 6817 6595 6851
rect 11253 6817 11287 6851
rect 14105 6817 14139 6851
rect 1409 6749 1443 6783
rect 2145 6749 2179 6783
rect 3801 6749 3835 6783
rect 4068 6749 4102 6783
rect 5641 6749 5675 6783
rect 7389 6749 7423 6783
rect 9873 6749 9907 6783
rect 10517 6749 10551 6783
rect 12081 6749 12115 6783
rect 12348 6749 12382 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 2053 6681 2087 6715
rect 2390 6681 2424 6715
rect 5917 6681 5951 6715
rect 7656 6681 7690 6715
rect 9045 6681 9079 6715
rect 9137 6681 9171 6715
rect 9689 6681 9723 6715
rect 10425 6681 10459 6715
rect 11345 6681 11379 6715
rect 11897 6681 11931 6715
rect 5181 6613 5215 6647
rect 7205 6613 7239 6647
rect 8769 6613 8803 6647
rect 10609 6613 10643 6647
rect 10793 6613 10827 6647
rect 3893 6409 3927 6443
rect 5549 6409 5583 6443
rect 6193 6409 6227 6443
rect 8309 6409 8343 6443
rect 8585 6409 8619 6443
rect 9045 6409 9079 6443
rect 14381 6409 14415 6443
rect 3157 6341 3191 6375
rect 4436 6341 4470 6375
rect 9505 6341 9539 6375
rect 10885 6341 10919 6375
rect 1409 6273 1443 6307
rect 1676 6273 1710 6307
rect 4077 6273 4111 6307
rect 5917 6273 5951 6307
rect 6009 6273 6043 6307
rect 7113 6273 7147 6307
rect 7573 6273 7607 6307
rect 8769 6273 8803 6307
rect 9229 6273 9263 6307
rect 10977 6273 11011 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12348 6273 12382 6307
rect 14197 6273 14231 6307
rect 14289 6273 14323 6307
rect 3065 6205 3099 6239
rect 4169 6205 4203 6239
rect 6469 6205 6503 6239
rect 7205 6205 7239 6239
rect 7665 6205 7699 6239
rect 7849 6205 7883 6239
rect 9413 6205 9447 6239
rect 10241 6205 10275 6239
rect 12081 6205 12115 6239
rect 13645 6205 13679 6239
rect 3617 6137 3651 6171
rect 5733 6137 5767 6171
rect 9965 6137 9999 6171
rect 11529 6137 11563 6171
rect 13461 6137 13495 6171
rect 2789 6069 2823 6103
rect 7021 6069 7055 6103
rect 7389 6069 7423 6103
rect 11069 6069 11103 6103
rect 11897 6069 11931 6103
rect 1593 5865 1627 5899
rect 3433 5865 3467 5899
rect 3985 5865 4019 5899
rect 4629 5865 4663 5899
rect 6469 5865 6503 5899
rect 7205 5865 7239 5899
rect 7573 5865 7607 5899
rect 8033 5865 8067 5899
rect 8401 5865 8435 5899
rect 11621 5865 11655 5899
rect 14105 5865 14139 5899
rect 3249 5797 3283 5831
rect 4813 5797 4847 5831
rect 10333 5797 10367 5831
rect 1869 5729 1903 5763
rect 2053 5729 2087 5763
rect 8953 5729 8987 5763
rect 10425 5729 10459 5763
rect 10609 5729 10643 5763
rect 11345 5729 11379 5763
rect 11897 5729 11931 5763
rect 13277 5729 13311 5763
rect 1777 5661 1811 5695
rect 3617 5661 3651 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 5356 5661 5390 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8309 5661 8343 5695
rect 8585 5661 8619 5695
rect 11161 5661 11195 5695
rect 12081 5661 12115 5695
rect 12725 5661 12759 5695
rect 14289 5661 14323 5695
rect 2513 5593 2547 5627
rect 2697 5593 2731 5627
rect 2789 5593 2823 5627
rect 9220 5593 9254 5627
rect 11069 5593 11103 5627
rect 13369 5593 13403 5627
rect 13921 5593 13955 5627
rect 4353 5525 4387 5559
rect 7757 5525 7791 5559
rect 8677 5525 8711 5559
rect 12541 5525 12575 5559
rect 12817 5525 12851 5559
rect 2237 5321 2271 5355
rect 5089 5321 5123 5355
rect 5825 5321 5859 5355
rect 6745 5321 6779 5355
rect 7389 5321 7423 5355
rect 11897 5321 11931 5355
rect 14289 5321 14323 5355
rect 2421 5253 2455 5287
rect 2605 5253 2639 5287
rect 6101 5253 6135 5287
rect 7849 5253 7883 5287
rect 10425 5253 10459 5287
rect 10517 5253 10551 5287
rect 13553 5253 13587 5287
rect 13645 5253 13679 5287
rect 2329 5185 2363 5219
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 6009 5185 6043 5219
rect 6561 5185 6595 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 7573 5185 7607 5219
rect 9689 5185 9723 5219
rect 9965 5185 9999 5219
rect 11345 5185 11379 5219
rect 11713 5185 11747 5219
rect 12256 5185 12290 5219
rect 14473 5185 14507 5219
rect 1685 5117 1719 5151
rect 4445 5117 4479 5151
rect 4629 5117 4663 5151
rect 5365 5117 5399 5151
rect 10701 5117 10735 5151
rect 11989 5117 12023 5151
rect 6837 5049 6871 5083
rect 9321 5049 9355 5083
rect 14105 5049 14139 5083
rect 7205 4981 7239 5015
rect 9781 4981 9815 5015
rect 10057 4981 10091 5015
rect 11161 4981 11195 5015
rect 13369 4981 13403 5015
rect 3249 4777 3283 4811
rect 4813 4777 4847 4811
rect 5549 4777 5583 4811
rect 10333 4777 10367 4811
rect 10885 4777 10919 4811
rect 11805 4777 11839 4811
rect 13369 4777 13403 4811
rect 3985 4709 4019 4743
rect 4169 4709 4203 4743
rect 9321 4709 9355 4743
rect 10517 4709 10551 4743
rect 12541 4709 12575 4743
rect 3065 4641 3099 4675
rect 6837 4641 6871 4675
rect 11989 4641 12023 4675
rect 12817 4641 12851 4675
rect 1409 4573 1443 4607
rect 2881 4573 2915 4607
rect 3801 4573 3835 4607
rect 4353 4573 4387 4607
rect 4445 4573 4479 4607
rect 4629 4573 4663 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 6009 4573 6043 4607
rect 6653 4573 6687 4607
rect 7389 4573 7423 4607
rect 8953 4573 8987 4607
rect 9137 4573 9171 4607
rect 9689 4573 9723 4607
rect 10425 4573 10459 4607
rect 11161 4573 11195 4607
rect 11345 4573 11379 4607
rect 14289 4573 14323 4607
rect 1676 4505 1710 4539
rect 7656 4505 7690 4539
rect 12081 4505 12115 4539
rect 13553 4505 13587 4539
rect 14381 4505 14415 4539
rect 2789 4437 2823 4471
rect 6561 4437 6595 4471
rect 7297 4437 7331 4471
rect 8769 4437 8803 4471
rect 13829 4437 13863 4471
rect 1777 4233 1811 4267
rect 3709 4233 3743 4267
rect 4445 4233 4479 4267
rect 5641 4233 5675 4267
rect 5733 4233 5767 4267
rect 7021 4233 7055 4267
rect 7481 4233 7515 4267
rect 8401 4233 8435 4267
rect 9137 4233 9171 4267
rect 14105 4165 14139 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 2145 4097 2179 4131
rect 2237 4097 2271 4131
rect 3065 4097 3099 4131
rect 3801 4097 3835 4131
rect 4905 4097 4939 4131
rect 5181 4097 5215 4131
rect 5917 4097 5951 4131
rect 6009 4097 6043 4131
rect 7389 4081 7423 4115
rect 7665 4097 7699 4131
rect 8677 4097 8711 4131
rect 9229 4097 9263 4131
rect 9689 4097 9723 4131
rect 9956 4097 9990 4131
rect 11345 4097 11379 4131
rect 12909 4097 12943 4131
rect 13185 4097 13219 4131
rect 13461 4097 13495 4131
rect 13921 4097 13955 4131
rect 2421 4029 2455 4063
rect 3249 4029 3283 4063
rect 3985 4029 4019 4063
rect 4997 4029 5031 4063
rect 6469 4029 6503 4063
rect 7849 4029 7883 4063
rect 8493 4029 8527 4063
rect 11529 4029 11563 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 13277 4029 13311 4063
rect 1501 3961 1535 3995
rect 4721 3961 4755 3995
rect 9321 3961 9355 3995
rect 11069 3961 11103 3995
rect 11161 3961 11195 3995
rect 1961 3893 1995 3927
rect 2605 3893 2639 3927
rect 6101 3893 6135 3927
rect 7205 3893 7239 3927
rect 12173 3893 12207 3927
rect 13001 3893 13035 3927
rect 14197 3893 14231 3927
rect 1777 3689 1811 3723
rect 2513 3689 2547 3723
rect 3617 3689 3651 3723
rect 4629 3689 4663 3723
rect 6285 3689 6319 3723
rect 7757 3689 7791 3723
rect 11437 3689 11471 3723
rect 11529 3689 11563 3723
rect 14289 3689 14323 3723
rect 4353 3621 4387 3655
rect 10701 3621 10735 3655
rect 13277 3621 13311 3655
rect 2053 3553 2087 3587
rect 2971 3553 3005 3587
rect 4077 3553 4111 3587
rect 8125 3553 8159 3587
rect 8401 3553 8435 3587
rect 8953 3553 8987 3587
rect 11897 3553 11931 3587
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 2697 3485 2731 3519
rect 3157 3485 3191 3519
rect 3893 3485 3927 3519
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 6377 3485 6411 3519
rect 9321 3485 9355 3519
rect 10793 3485 10827 3519
rect 11713 3485 11747 3519
rect 13461 3485 13495 3519
rect 14105 3485 14139 3519
rect 5172 3417 5206 3451
rect 6644 3417 6678 3451
rect 8217 3417 8251 3451
rect 9588 3417 9622 3451
rect 12142 3417 12176 3451
rect 13829 3417 13863 3451
rect 2789 3349 2823 3383
rect 2145 3145 2179 3179
rect 3249 3145 3283 3179
rect 3433 3145 3467 3179
rect 4261 3145 4295 3179
rect 4445 3145 4479 3179
rect 7021 3145 7055 3179
rect 9505 3145 9539 3179
rect 11253 3145 11287 3179
rect 12173 3145 12207 3179
rect 7297 3077 7331 3111
rect 7849 3077 7883 3111
rect 8585 3077 8619 3111
rect 8769 3077 8803 3111
rect 8861 3077 8895 3111
rect 10140 3077 10174 3111
rect 12357 3077 12391 3111
rect 12449 3077 12483 3111
rect 13001 3077 13035 3111
rect 1409 3009 1443 3043
rect 1685 3009 1719 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 4353 3009 4387 3043
rect 4813 3009 4847 3043
rect 4997 3009 5031 3043
rect 6469 3009 6503 3043
rect 7941 3009 7975 3043
rect 9689 3009 9723 3043
rect 11621 3009 11655 3043
rect 13185 3009 13219 3043
rect 13645 3009 13679 3043
rect 3801 2941 3835 2975
rect 5549 2941 5583 2975
rect 5733 2941 5767 2975
rect 7205 2941 7239 2975
rect 8125 2941 8159 2975
rect 9045 2941 9079 2975
rect 9873 2941 9907 2975
rect 13921 2941 13955 2975
rect 1501 2873 1535 2907
rect 6193 2873 6227 2907
rect 1869 2805 1903 2839
rect 2421 2805 2455 2839
rect 5457 2805 5491 2839
rect 13277 2805 13311 2839
rect 2789 2601 2823 2635
rect 4445 2601 4479 2635
rect 5549 2601 5583 2635
rect 9781 2601 9815 2635
rect 11345 2601 11379 2635
rect 14105 2601 14139 2635
rect 2421 2533 2455 2567
rect 3617 2533 3651 2567
rect 4169 2533 4203 2567
rect 4997 2533 5031 2567
rect 10609 2533 10643 2567
rect 13001 2533 13035 2567
rect 13829 2533 13863 2567
rect 1409 2465 1443 2499
rect 5181 2465 5215 2499
rect 7021 2465 7055 2499
rect 7665 2465 7699 2499
rect 10701 2465 10735 2499
rect 10885 2465 10919 2499
rect 11897 2465 11931 2499
rect 13277 2465 13311 2499
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 3157 2397 3191 2431
rect 3433 2397 3467 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 4353 2397 4387 2431
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 5365 2397 5399 2431
rect 6469 2397 6503 2431
rect 7849 2397 7883 2431
rect 8217 2397 8251 2431
rect 8401 2397 8435 2431
rect 9045 2397 9079 2431
rect 9689 2397 9723 2431
rect 10057 2397 10091 2431
rect 14289 2397 14323 2431
rect 6009 2329 6043 2363
rect 7113 2329 7147 2363
rect 8769 2329 8803 2363
rect 11621 2329 11655 2363
rect 11713 2329 11747 2363
rect 12449 2329 12483 2363
rect 12541 2329 12575 2363
rect 13369 2329 13403 2363
rect 2973 2261 3007 2295
rect 3341 2261 3375 2295
rect 3985 2261 4019 2295
rect 4721 2261 4755 2295
rect 6745 2261 6779 2295
rect 9137 2261 9171 2295
<< metal1 >>
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13780 17292 13829 17320
rect 13780 17280 13786 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 2774 17212 2780 17264
rect 2832 17212 2838 17264
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 1872 17116 1900 17147
rect 2406 17144 2412 17196
rect 2464 17144 2470 17196
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 11020 17156 13553 17184
rect 11020 17144 11026 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 14568 17184 14596 17280
rect 14507 17156 14596 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 5626 17116 5632 17128
rect 1872 17088 5632 17116
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 1026 16940 1032 16992
rect 1084 16980 1090 16992
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1084 16952 1961 16980
rect 1084 16940 1090 16952
rect 1949 16949 1961 16952
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 14274 16940 14280 16992
rect 14332 16940 14338 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 934 16736 940 16788
rect 992 16776 998 16788
rect 1765 16779 1823 16785
rect 1765 16776 1777 16779
rect 992 16748 1777 16776
rect 992 16736 998 16748
rect 1765 16745 1777 16748
rect 1811 16745 1823 16779
rect 1765 16739 1823 16745
rect 2225 16779 2283 16785
rect 2225 16745 2237 16779
rect 2271 16776 2283 16779
rect 2406 16776 2412 16788
rect 2271 16748 2412 16776
rect 2271 16745 2283 16748
rect 2225 16739 2283 16745
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 14642 16736 14648 16788
rect 14700 16736 14706 16788
rect 9858 16640 9864 16652
rect 2148 16612 9864 16640
rect 2148 16581 2176 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 14660 16640 14688 16736
rect 13924 16612 14688 16640
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 8754 16572 8760 16584
rect 8435 16544 8760 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 13924 16581 13952 16612
rect 13909 16575 13967 16581
rect 13909 16541 13921 16575
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 15010 16572 15016 16584
rect 14323 16544 15016 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 1673 16507 1731 16513
rect 1673 16473 1685 16507
rect 1719 16504 1731 16507
rect 1719 16476 2774 16504
rect 1719 16473 1731 16476
rect 1673 16467 1731 16473
rect 2746 16436 2774 16476
rect 8205 16439 8263 16445
rect 8205 16436 8217 16439
rect 2746 16408 8217 16436
rect 8205 16405 8217 16408
rect 8251 16405 8263 16439
rect 8205 16399 8263 16405
rect 13722 16396 13728 16448
rect 13780 16396 13786 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14461 16439 14519 16445
rect 14461 16436 14473 16439
rect 13872 16408 14473 16436
rect 13872 16396 13878 16408
rect 14461 16405 14473 16408
rect 14507 16405 14519 16439
rect 14461 16399 14519 16405
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 934 16192 940 16244
rect 992 16232 998 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 992 16204 1593 16232
rect 992 16192 998 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 9950 16096 9956 16108
rect 1535 16068 9956 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 1176 15660 2145 15688
rect 1176 15648 1182 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 13814 15688 13820 15700
rect 2133 15651 2191 15657
rect 12406 15660 13820 15688
rect 1489 15487 1547 15493
rect 1489 15453 1501 15487
rect 1535 15484 1547 15487
rect 3418 15484 3424 15496
rect 1535 15456 3424 15484
rect 1535 15453 1547 15456
rect 1489 15447 1547 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 12406 15484 12434 15660
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 14415 15660 14872 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 14844 15632 14872 15660
rect 14826 15580 14832 15632
rect 14884 15580 14890 15632
rect 5675 15456 12434 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 13964 15456 14197 15484
rect 13964 15444 13970 15456
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 2041 15419 2099 15425
rect 2041 15385 2053 15419
rect 2087 15416 2099 15419
rect 2866 15416 2872 15428
rect 2087 15388 2872 15416
rect 2087 15385 2099 15388
rect 2041 15379 2099 15385
rect 2866 15376 2872 15388
rect 2924 15376 2930 15428
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 5902 15348 5908 15360
rect 5767 15320 5908 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 8202 15144 8208 15156
rect 2516 15116 8208 15144
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 1670 15008 1676 15020
rect 1627 14980 1676 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2516 15017 2544 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 2593 15079 2651 15085
rect 2593 15045 2605 15079
rect 2639 15076 2651 15079
rect 7190 15076 7196 15088
rect 2639 15048 7196 15076
rect 2639 15045 2651 15048
rect 2593 15039 2651 15045
rect 7190 15036 7196 15048
rect 7248 15036 7254 15088
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 12066 15076 12072 15088
rect 10008 15048 12072 15076
rect 10008 15036 10014 15048
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 1964 14980 2237 15008
rect 1964 14816 1992 14980
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 2792 14940 2820 14971
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 4890 15008 4896 15020
rect 3099 14980 4896 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 10836 14980 14197 15008
rect 10836 14968 10842 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 4154 14940 4160 14952
rect 2792 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 2409 14875 2467 14881
rect 2409 14841 2421 14875
rect 2455 14872 2467 14875
rect 3602 14872 3608 14884
rect 2455 14844 3608 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 3602 14832 3608 14844
rect 3660 14832 3666 14884
rect 1394 14764 1400 14816
rect 1452 14764 1458 14816
rect 1946 14764 1952 14816
rect 2004 14764 2010 14816
rect 3234 14764 3240 14816
rect 3292 14764 3298 14816
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 9122 14804 9128 14816
rect 3384 14776 9128 14804
rect 3384 14764 3390 14776
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1452 14572 3372 14600
rect 1452 14560 1458 14572
rect 1765 14535 1823 14541
rect 1765 14501 1777 14535
rect 1811 14501 1823 14535
rect 1765 14495 1823 14501
rect 1780 14464 1808 14495
rect 1780 14436 2360 14464
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 2332 14405 2360 14436
rect 2406 14424 2412 14476
rect 2464 14424 2470 14476
rect 3344 14464 3372 14572
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 10226 14600 10232 14612
rect 3568 14572 10232 14600
rect 3568 14560 3574 14572
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9916 14504 10057 14532
rect 9916 14492 9922 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 3344 14436 3464 14464
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1912 14368 1961 14396
rect 1912 14356 1918 14368
rect 1949 14365 1961 14368
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 2958 14396 2964 14408
rect 2915 14368 2964 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 2240 14328 2268 14359
rect 2958 14356 2964 14368
rect 3016 14396 3022 14408
rect 3436 14405 3464 14436
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 9950 14464 9956 14476
rect 3752 14436 9956 14464
rect 3752 14424 3758 14436
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 3016 14368 3157 14396
rect 3016 14356 3022 14368
rect 3145 14365 3157 14368
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3510 14356 3516 14408
rect 3568 14356 3574 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8352 14368 8585 14396
rect 8352 14356 8358 14368
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 10689 14399 10747 14405
rect 10459 14368 10548 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 3528 14328 3556 14356
rect 2240 14300 3556 14328
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 9306 14328 9312 14340
rect 3844 14300 9312 14328
rect 3844 14288 3850 14300
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9490 14288 9496 14340
rect 9548 14288 9554 14340
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14297 9643 14331
rect 9585 14291 9643 14297
rect 1673 14263 1731 14269
rect 1673 14229 1685 14263
rect 1719 14260 1731 14263
rect 1854 14260 1860 14272
rect 1719 14232 1860 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2038 14220 2044 14272
rect 2096 14220 2102 14272
rect 3326 14220 3332 14272
rect 3384 14220 3390 14272
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3605 14263 3663 14269
rect 3605 14260 3617 14263
rect 3568 14232 3617 14260
rect 3568 14220 3574 14232
rect 3605 14229 3617 14232
rect 3651 14229 3663 14263
rect 3605 14223 3663 14229
rect 4065 14263 4123 14269
rect 4065 14229 4077 14263
rect 4111 14260 4123 14263
rect 5258 14260 5264 14272
rect 4111 14232 5264 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 8386 14220 8392 14272
rect 8444 14220 8450 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8536 14232 8953 14260
rect 8536 14220 8542 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 9600 14260 9628 14291
rect 10520 14269 10548 14368
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10962 14396 10968 14408
rect 10735 14368 10968 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 10229 14263 10287 14269
rect 10229 14260 10241 14263
rect 9600 14232 10241 14260
rect 8941 14223 8999 14229
rect 10229 14229 10241 14232
rect 10275 14229 10287 14263
rect 10229 14223 10287 14229
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14229 10563 14263
rect 10505 14223 10563 14229
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1210 14016 1216 14068
rect 1268 14056 1274 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 1268 14028 2881 14056
rect 1268 14016 1274 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 3050 14016 3056 14068
rect 3108 14016 3114 14068
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 3694 14056 3700 14068
rect 3528 14028 3700 14056
rect 1486 13948 1492 14000
rect 1544 13948 1550 14000
rect 1670 13948 1676 14000
rect 1728 13988 1734 14000
rect 2777 13991 2835 13997
rect 1728 13960 2268 13988
rect 1728 13948 1734 13960
rect 474 13880 480 13932
rect 532 13920 538 13932
rect 2240 13929 2268 13960
rect 2777 13957 2789 13991
rect 2823 13988 2835 13991
rect 3068 13988 3096 14016
rect 2823 13960 3372 13988
rect 2823 13957 2835 13960
rect 2777 13951 2835 13957
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 532 13892 1961 13920
rect 532 13880 538 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 2314 13880 2320 13932
rect 2372 13880 2378 13932
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 3344 13929 3372 13960
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2556 13892 3065 13920
rect 2556 13880 2562 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 3528 13852 3556 14028
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 5074 14056 5080 14068
rect 3927 14028 5080 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 8570 14016 8576 14068
rect 8628 14056 8634 14068
rect 9490 14056 9496 14068
rect 8628 14028 9496 14056
rect 8628 14016 8634 14028
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 10962 14016 10968 14068
rect 11020 14016 11026 14068
rect 13722 14016 13728 14068
rect 13780 14016 13786 14068
rect 3786 13988 3792 14000
rect 3620 13960 3792 13988
rect 3620 13929 3648 13960
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 4798 13988 4804 14000
rect 3988 13960 4804 13988
rect 3988 13929 4016 13960
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 9677 13991 9735 13997
rect 9677 13957 9689 13991
rect 9723 13988 9735 13991
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 9723 13960 10425 13988
rect 9723 13957 9735 13960
rect 9677 13951 9735 13957
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10413 13951 10471 13957
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 3712 13852 3740 13883
rect 4062 13880 4068 13932
rect 4120 13880 4126 13932
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 2087 13824 3556 13852
rect 3620 13824 3740 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 750 13744 756 13796
rect 808 13784 814 13796
rect 3418 13784 3424 13796
rect 808 13756 3424 13784
rect 808 13744 814 13756
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 3510 13744 3516 13796
rect 3568 13784 3574 13796
rect 3620 13784 3648 13824
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 4448 13852 4476 13883
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 10980 13920 11008 14016
rect 10376 13892 11008 13920
rect 12621 13923 12679 13929
rect 10376 13880 10382 13892
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13740 13920 13768 14016
rect 12667 13892 13768 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 6914 13852 6920 13864
rect 3844 13824 4476 13852
rect 4540 13824 6920 13852
rect 3844 13812 3850 13824
rect 3568 13756 3648 13784
rect 4249 13787 4307 13793
rect 3568 13744 3574 13756
rect 4249 13753 4261 13787
rect 4295 13784 4307 13787
rect 4540 13784 4568 13824
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 7708 13824 7941 13852
rect 7708 13812 7714 13824
rect 7929 13821 7941 13824
rect 7975 13821 7987 13855
rect 7929 13815 7987 13821
rect 8110 13812 8116 13864
rect 8168 13812 8174 13864
rect 8662 13812 8668 13864
rect 8720 13812 8726 13864
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9272 13824 9597 13852
rect 9272 13812 9278 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14458 13852 14464 13864
rect 14415 13824 14464 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 10870 13784 10876 13796
rect 4295 13756 4568 13784
rect 9232 13756 10876 13784
rect 4295 13753 4307 13756
rect 4249 13747 4307 13753
rect 1578 13676 1584 13728
rect 1636 13676 1642 13728
rect 3145 13719 3203 13725
rect 3145 13685 3157 13719
rect 3191 13716 3203 13719
rect 3234 13716 3240 13728
rect 3191 13688 3240 13716
rect 3191 13685 3203 13688
rect 3145 13679 3203 13685
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 9232 13716 9260 13756
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 3384 13688 9260 13716
rect 3384 13676 3390 13688
rect 9306 13676 9312 13728
rect 9364 13676 9370 13728
rect 12710 13676 12716 13728
rect 12768 13676 12774 13728
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 3053 13515 3111 13521
rect 3053 13481 3065 13515
rect 3099 13512 3111 13515
rect 7745 13515 7803 13521
rect 3099 13484 7328 13512
rect 3099 13481 3111 13484
rect 3053 13475 3111 13481
rect 1118 13404 1124 13456
rect 1176 13444 1182 13456
rect 1176 13416 2912 13444
rect 1176 13404 1182 13416
rect 566 13336 572 13388
rect 624 13376 630 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 624 13348 2513 13376
rect 624 13336 630 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 2130 13268 2136 13320
rect 2188 13268 2194 13320
rect 2884 13317 2912 13416
rect 3234 13336 3240 13388
rect 3292 13376 3298 13388
rect 3292 13348 5120 13376
rect 3292 13336 3298 13348
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3326 13308 3332 13320
rect 3191 13280 3332 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 658 13200 664 13252
rect 716 13240 722 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 716 13212 1501 13240
rect 716 13200 722 13212
rect 1489 13209 1501 13212
rect 1535 13209 1547 13243
rect 2424 13240 2452 13271
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 5092 13317 5120 13348
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 2958 13240 2964 13252
rect 2424 13212 2964 13240
rect 1489 13203 1547 13209
rect 2958 13200 2964 13212
rect 3016 13200 3022 13252
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 992 13144 1593 13172
rect 992 13132 998 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 2314 13132 2320 13184
rect 2372 13132 2378 13184
rect 3326 13132 3332 13184
rect 3384 13132 3390 13184
rect 3602 13132 3608 13184
rect 3660 13132 3666 13184
rect 3804 13172 3832 13271
rect 4080 13240 4108 13271
rect 5994 13240 6000 13252
rect 4080 13212 6000 13240
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 4982 13172 4988 13184
rect 3804 13144 4988 13172
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5166 13132 5172 13184
rect 5224 13132 5230 13184
rect 7300 13172 7328 13484
rect 7745 13481 7757 13515
rect 7791 13512 7803 13515
rect 8110 13512 8116 13524
rect 7791 13484 8116 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8294 13472 8300 13524
rect 8352 13472 8358 13524
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8812 13484 10272 13512
rect 8812 13472 8818 13484
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13444 7435 13447
rect 8312 13444 8340 13472
rect 7423 13416 8340 13444
rect 10244 13444 10272 13484
rect 10318 13472 10324 13524
rect 10376 13472 10382 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 10428 13484 13921 13512
rect 10428 13444 10456 13484
rect 13909 13481 13921 13484
rect 13955 13481 13967 13515
rect 13909 13475 13967 13481
rect 14274 13472 14280 13524
rect 14332 13472 14338 13524
rect 14292 13444 14320 13472
rect 10244 13416 10456 13444
rect 12406 13416 14320 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8386 13376 8392 13388
rect 8159 13348 8392 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7607 13280 7665 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13308 7987 13311
rect 8478 13308 8484 13320
rect 7975 13280 8484 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 7668 13240 7696 13271
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13308 8999 13311
rect 11054 13308 11060 13320
rect 8987 13280 11060 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 11054 13268 11060 13280
rect 11112 13308 11118 13320
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 11112 13280 11253 13308
rect 11112 13268 11118 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11508 13311 11566 13317
rect 11508 13277 11520 13311
rect 11554 13308 11566 13311
rect 12406 13308 12434 13416
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12768 13348 12817 13376
rect 12768 13336 12774 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 11554 13280 12434 13308
rect 11554 13277 11566 13280
rect 11508 13271 11566 13277
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 8386 13240 8392 13252
rect 7668 13212 8392 13240
rect 8386 13200 8392 13212
rect 8444 13240 8450 13252
rect 8662 13240 8668 13252
rect 8444 13212 8668 13240
rect 8444 13200 8450 13212
rect 8662 13200 8668 13212
rect 8720 13200 8726 13252
rect 9208 13243 9266 13249
rect 9208 13209 9220 13243
rect 9254 13240 9266 13243
rect 9306 13240 9312 13252
rect 9254 13212 9312 13240
rect 9254 13209 9266 13212
rect 9208 13203 9266 13209
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 13740 13240 13768 13271
rect 14182 13268 14188 13320
rect 14240 13268 14246 13320
rect 12308 13212 13768 13240
rect 12308 13200 12314 13212
rect 11606 13172 11612 13184
rect 7300 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 12618 13132 12624 13184
rect 12676 13132 12682 13184
rect 13446 13132 13452 13184
rect 13504 13132 13510 13184
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 2188 12940 3525 12968
rect 2188 12928 2194 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 8297 12971 8355 12977
rect 3513 12931 3571 12937
rect 3896 12940 5028 12968
rect 382 12860 388 12912
rect 440 12900 446 12912
rect 3896 12900 3924 12940
rect 440 12872 3924 12900
rect 3973 12903 4031 12909
rect 440 12860 446 12872
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 4246 12900 4252 12912
rect 4019 12872 4252 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 4522 12860 4528 12912
rect 4580 12900 4586 12912
rect 5000 12909 5028 12940
rect 8297 12937 8309 12971
rect 8343 12968 8355 12971
rect 8343 12940 8524 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 4985 12903 5043 12909
rect 4580 12872 4752 12900
rect 4580 12860 4586 12872
rect 1762 12792 1768 12844
rect 1820 12792 1826 12844
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2038 12832 2044 12844
rect 1903 12804 2044 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 860 12736 2329 12764
rect 860 12640 888 12736
rect 2317 12733 2329 12736
rect 2363 12764 2375 12767
rect 2884 12764 2912 12795
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3016 12804 3709 12832
rect 3016 12792 3022 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2363 12736 2912 12764
rect 2976 12736 3065 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2976 12708 3004 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 1995 12668 2912 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 842 12588 848 12640
rect 900 12588 906 12640
rect 1578 12588 1584 12640
rect 1636 12588 1642 12640
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2464 12600 2697 12628
rect 2464 12588 2470 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2884 12628 2912 12668
rect 2958 12656 2964 12708
rect 3016 12656 3022 12708
rect 3712 12696 3740 12795
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 4724 12841 4752 12872
rect 4985 12869 4997 12903
rect 5031 12869 5043 12903
rect 4985 12863 5043 12869
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 7098 12900 7104 12912
rect 5583 12872 7104 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 8496 12900 8524 12940
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 11790 12968 11796 12980
rect 8628 12940 11796 12968
rect 8628 12928 8634 12940
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12345 12971 12403 12977
rect 12345 12937 12357 12971
rect 12391 12968 12403 12971
rect 12986 12968 12992 12980
rect 12391 12940 12992 12968
rect 12391 12937 12403 12940
rect 12345 12931 12403 12937
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13541 12971 13599 12977
rect 13541 12968 13553 12971
rect 13372 12940 13553 12968
rect 11514 12900 11520 12912
rect 8496 12872 9536 12900
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5491 12804 5672 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4062 12764 4068 12776
rect 3927 12736 4068 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4908 12764 4936 12795
rect 5258 12764 5264 12776
rect 4396 12736 5264 12764
rect 4396 12724 4402 12736
rect 5258 12724 5264 12736
rect 5316 12764 5322 12776
rect 5368 12764 5396 12795
rect 5316 12736 5396 12764
rect 5316 12724 5322 12736
rect 5644 12696 5672 12804
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 7000 12835 7058 12841
rect 7000 12801 7012 12835
rect 7046 12832 7058 12835
rect 7282 12832 7288 12844
rect 7046 12804 7288 12832
rect 7046 12801 7058 12804
rect 7000 12795 7058 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 8527 12804 8708 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 5810 12724 5816 12776
rect 5868 12724 5874 12776
rect 6730 12724 6736 12776
rect 6788 12724 6794 12776
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8352 12736 8585 12764
rect 8352 12724 8358 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 8113 12699 8171 12705
rect 3712 12668 5580 12696
rect 5644 12668 6776 12696
rect 3234 12628 3240 12640
rect 2884 12600 3240 12628
rect 2685 12591 2743 12597
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 5552 12628 5580 12668
rect 6638 12628 6644 12640
rect 5552 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 6748 12628 6776 12668
rect 8113 12665 8125 12699
rect 8159 12696 8171 12699
rect 8386 12696 8392 12708
rect 8159 12668 8392 12696
rect 8159 12665 8171 12668
rect 8113 12659 8171 12665
rect 8386 12656 8392 12668
rect 8444 12696 8450 12708
rect 8680 12696 8708 12804
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9508 12841 9536 12872
rect 11072 12872 11520 12900
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10410 12832 10416 12844
rect 10367 12804 10416 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10410 12792 10416 12804
rect 10468 12832 10474 12844
rect 11072 12841 11100 12872
rect 11514 12860 11520 12872
rect 11572 12900 11578 12912
rect 11572 12872 12296 12900
rect 11572 12860 11578 12872
rect 12268 12841 12296 12872
rect 12618 12860 12624 12912
rect 12676 12860 12682 12912
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10468 12804 11069 12832
rect 10468 12792 10474 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12636 12832 12664 12860
rect 12299 12804 12664 12832
rect 12989 12835 13047 12841
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 13372 12832 13400 12940
rect 13541 12937 13553 12940
rect 13587 12937 13599 12971
rect 13541 12931 13599 12937
rect 13924 12872 14136 12900
rect 13311 12804 13400 12832
rect 13725 12835 13783 12841
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13924 12832 13952 12872
rect 14108 12841 14136 12872
rect 13771 12804 13952 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 8757 12767 8815 12773
rect 8757 12733 8769 12767
rect 8803 12764 8815 12767
rect 11348 12764 11376 12795
rect 8803 12736 9352 12764
rect 8803 12733 8815 12736
rect 8757 12727 8815 12733
rect 9030 12696 9036 12708
rect 8444 12668 9036 12696
rect 8444 12656 8450 12668
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 9324 12705 9352 12736
rect 10888 12736 11376 12764
rect 13004 12764 13032 12795
rect 13004 12736 13860 12764
rect 10888 12705 10916 12736
rect 9309 12699 9367 12705
rect 9309 12665 9321 12699
rect 9355 12665 9367 12699
rect 9309 12659 9367 12665
rect 10873 12699 10931 12705
rect 10873 12665 10885 12699
rect 10919 12665 10931 12699
rect 10873 12659 10931 12665
rect 11164 12668 12434 12696
rect 8662 12628 8668 12640
rect 6748 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 11164 12637 11192 12668
rect 12406 12640 12434 12668
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 13832 12705 13860 12736
rect 13817 12699 13875 12705
rect 12768 12668 13676 12696
rect 12768 12656 12774 12668
rect 11149 12631 11207 12637
rect 11149 12597 11161 12631
rect 11195 12597 11207 12631
rect 12406 12600 12440 12640
rect 11149 12591 11207 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 13173 12631 13231 12637
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 13262 12628 13268 12640
rect 13219 12600 13268 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 13449 12631 13507 12637
rect 13449 12597 13461 12631
rect 13495 12628 13507 12631
rect 13538 12628 13544 12640
rect 13495 12600 13544 12628
rect 13495 12597 13507 12600
rect 13449 12591 13507 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13648 12628 13676 12668
rect 13817 12665 13829 12699
rect 13863 12665 13875 12699
rect 13817 12659 13875 12665
rect 13924 12628 13952 12804
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14016 12764 14044 12795
rect 14458 12764 14464 12776
rect 14016 12736 14464 12764
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 13648 12600 13952 12628
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14550 12628 14556 12640
rect 14231 12600 14556 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 2593 12427 2651 12433
rect 2593 12424 2605 12427
rect 2556 12396 2605 12424
rect 2556 12384 2562 12396
rect 2593 12393 2605 12396
rect 2639 12393 2651 12427
rect 2593 12387 2651 12393
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 4062 12424 4068 12436
rect 3476 12396 4068 12424
rect 3476 12384 3482 12396
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 7282 12384 7288 12436
rect 7340 12384 7346 12436
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 7423 12396 7880 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 2424 12328 4016 12356
rect 2424 12229 2452 12328
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 3878 12288 3884 12300
rect 3568 12260 3884 12288
rect 3568 12248 3574 12260
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 3988 12288 4016 12328
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 6273 12359 6331 12365
rect 4212 12328 4476 12356
rect 4212 12316 4218 12328
rect 4338 12288 4344 12300
rect 3988 12260 4344 12288
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4448 12297 4476 12328
rect 6273 12325 6285 12359
rect 6319 12356 6331 12359
rect 6319 12328 6868 12356
rect 6319 12325 6331 12328
rect 6273 12319 6331 12325
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 6730 12288 6736 12300
rect 4433 12251 4491 12257
rect 5920 12260 6736 12288
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2961 12223 3019 12229
rect 2961 12220 2973 12223
rect 2731 12192 2973 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2961 12189 2973 12192
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5534 12220 5540 12232
rect 4939 12192 5540 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 1486 12112 1492 12164
rect 1544 12112 1550 12164
rect 2148 12152 2176 12183
rect 2498 12152 2504 12164
rect 2148 12124 2504 12152
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 3160 12152 3188 12183
rect 2924 12124 3188 12152
rect 2924 12112 2930 12124
rect 934 12044 940 12096
rect 992 12084 998 12096
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 992 12056 1593 12084
rect 992 12044 998 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 3234 12084 3240 12096
rect 1995 12056 3240 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3602 12084 3608 12096
rect 3476 12056 3608 12084
rect 3476 12044 3482 12056
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3786 12044 3792 12096
rect 3844 12044 3850 12096
rect 3988 12084 4016 12183
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 5920 12220 5948 12260
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 6840 12232 6868 12328
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7852 12297 7880 12396
rect 9214 12384 9220 12436
rect 9272 12424 9278 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 9272 12396 9321 12424
rect 9272 12384 9278 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 12897 12427 12955 12433
rect 12897 12393 12909 12427
rect 12943 12424 12955 12427
rect 12986 12424 12992 12436
rect 12943 12396 12992 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 12986 12384 12992 12396
rect 13044 12424 13050 12436
rect 13446 12424 13452 12436
rect 13044 12396 13452 12424
rect 13044 12384 13050 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14182 12424 14188 12436
rect 13771 12396 14188 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 10689 12359 10747 12365
rect 7944 12328 9904 12356
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7248 12260 7665 12288
rect 7248 12248 7254 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 5592 12192 5948 12220
rect 5592 12180 5598 12192
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 6052 12192 6377 12220
rect 6052 12180 6058 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6822 12220 6828 12232
rect 6687 12192 6828 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7668 12220 7696 12251
rect 7944 12220 7972 12328
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12288 9183 12291
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 9171 12260 9781 12288
rect 9171 12257 9183 12260
rect 9125 12251 9183 12257
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 9876 12288 9904 12328
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 11149 12359 11207 12365
rect 11149 12356 11161 12359
rect 10735 12328 11161 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 11149 12325 11161 12328
rect 11195 12356 11207 12359
rect 11195 12328 13032 12356
rect 11195 12325 11207 12328
rect 11149 12319 11207 12325
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 9876 12260 10793 12288
rect 9769 12251 9827 12257
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 12158 12248 12164 12300
rect 12216 12248 12222 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 13004 12297 13032 12328
rect 14366 12316 14372 12368
rect 14424 12316 14430 12368
rect 12989 12291 13047 12297
rect 12989 12257 13001 12291
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7668 12192 7972 12220
rect 8036 12192 8401 12220
rect 4154 12112 4160 12164
rect 4212 12112 4218 12164
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12152 4307 12155
rect 4522 12152 4528 12164
rect 4295 12124 4528 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 5160 12155 5218 12161
rect 5160 12121 5172 12155
rect 5206 12152 5218 12155
rect 5350 12152 5356 12164
rect 5206 12124 5356 12152
rect 5206 12121 5218 12124
rect 5160 12115 5218 12121
rect 5350 12112 5356 12124
rect 5408 12112 5414 12164
rect 4706 12084 4712 12096
rect 3988 12056 4712 12084
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 5684 12056 6469 12084
rect 5684 12044 5690 12056
rect 6457 12053 6469 12056
rect 6503 12053 6515 12087
rect 6840 12084 6868 12180
rect 8036 12084 8064 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9088 12192 9689 12220
rect 9088 12180 9094 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 8496 12152 8524 12180
rect 10060 12152 10088 12183
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 11204 12192 12265 12220
rect 11204 12180 11210 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 13170 12180 13176 12232
rect 13228 12180 13234 12232
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12189 13967 12223
rect 13909 12183 13967 12189
rect 8496 12124 10088 12152
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12342 12152 12348 12164
rect 11664 12124 12348 12152
rect 11664 12112 11670 12124
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 13924 12152 13952 12183
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 12452 12124 13952 12152
rect 6840 12056 8064 12084
rect 6457 12047 6515 12053
rect 8294 12044 8300 12096
rect 8352 12044 8358 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 12452 12084 12480 12124
rect 10100 12056 12480 12084
rect 10100 12044 10106 12056
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1544 11852 2145 11880
rect 1544 11840 1550 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2866 11880 2872 11892
rect 2639 11852 2872 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 2976 11852 3556 11880
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 2976 11812 3004 11852
rect 3418 11812 3424 11824
rect 1903 11784 3004 11812
rect 3068 11784 3424 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11744 1455 11747
rect 1670 11744 1676 11756
rect 1443 11716 1676 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 1780 11676 1808 11707
rect 2038 11704 2044 11756
rect 2096 11704 2102 11756
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2777 11747 2835 11753
rect 2363 11716 2544 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2406 11676 2412 11688
rect 1780 11648 2412 11676
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 1210 11568 1216 11620
rect 1268 11608 1274 11620
rect 1268 11580 2452 11608
rect 1268 11568 1274 11580
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 1489 11543 1547 11549
rect 1489 11540 1501 11543
rect 1452 11512 1501 11540
rect 1452 11500 1458 11512
rect 1489 11509 1501 11512
rect 1535 11509 1547 11543
rect 1489 11503 1547 11509
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 2130 11540 2136 11552
rect 1728 11512 2136 11540
rect 1728 11500 1734 11512
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2424 11549 2452 11580
rect 2516 11552 2544 11716
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 3068 11744 3096 11784
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 3528 11812 3556 11852
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 3844 11852 4200 11880
rect 3844 11840 3850 11852
rect 3528 11784 4108 11812
rect 3142 11753 3148 11756
rect 2823 11716 3096 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 3136 11707 3148 11753
rect 3142 11704 3148 11707
rect 3200 11704 3206 11756
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11645 2927 11679
rect 4080 11676 4108 11784
rect 4172 11744 4200 11852
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4304 11852 4445 11880
rect 4304 11840 4310 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 5350 11840 5356 11892
rect 5408 11840 5414 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7558 11880 7564 11892
rect 7147 11852 7564 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 8294 11840 8300 11892
rect 8352 11840 8358 11892
rect 8478 11840 8484 11892
rect 8536 11840 8542 11892
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10226 11880 10232 11892
rect 9999 11852 10232 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 10962 11880 10968 11892
rect 10367 11852 10968 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11146 11840 11152 11892
rect 11204 11840 11210 11892
rect 11977 11883 12035 11889
rect 11977 11849 11989 11883
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 13170 11880 13176 11892
rect 12299 11852 13176 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 6880 11784 7328 11812
rect 6880 11772 6886 11784
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4172 11716 4629 11744
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 7300 11753 7328 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8386 11812 8392 11824
rect 7708 11784 8392 11812
rect 7708 11772 7714 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6052 11716 7021 11744
rect 6052 11704 6058 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7466 11744 7472 11756
rect 7331 11716 7472 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 8496 11744 8524 11840
rect 10410 11772 10416 11824
rect 10468 11772 10474 11824
rect 7883 11716 8524 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 4080 11648 4844 11676
rect 2869 11639 2927 11645
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 2498 11500 2504 11552
rect 2556 11500 2562 11552
rect 2884 11540 2912 11639
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 4706 11608 4712 11620
rect 4295 11580 4712 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 4816 11608 4844 11648
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 5224 11648 5457 11676
rect 5224 11636 5230 11648
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7576 11676 7604 11707
rect 10134 11704 10140 11756
rect 10192 11704 10198 11756
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10428 11744 10456 11772
rect 10275 11716 10456 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 6972 11648 7604 11676
rect 7653 11679 7711 11685
rect 6972 11636 6978 11648
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 11164 11676 11192 11840
rect 11992 11812 12020 11843
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13630 11840 13636 11892
rect 13688 11840 13694 11892
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14182 11880 14188 11892
rect 14047 11852 14188 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 7699 11648 11192 11676
rect 11808 11784 12020 11812
rect 12176 11784 12572 11812
rect 11808 11676 11836 11784
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12176 11753 12204 11784
rect 12544 11753 12572 11784
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11940 11716 12173 11744
rect 11940 11704 11946 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12667 11716 13185 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 12452 11676 12480 11707
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13320 11716 13921 11744
rect 13320 11704 13326 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 11808 11648 12480 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 4816 11580 6224 11608
rect 3970 11540 3976 11552
rect 2884 11512 3976 11540
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 6089 11543 6147 11549
rect 6089 11540 6101 11543
rect 5776 11512 6101 11540
rect 5776 11500 5782 11512
rect 6089 11509 6101 11512
rect 6135 11509 6147 11543
rect 6196 11540 6224 11580
rect 6822 11568 6828 11620
rect 6880 11568 6886 11620
rect 7668 11608 7696 11639
rect 12986 11636 12992 11688
rect 13044 11636 13050 11688
rect 6932 11580 7696 11608
rect 11716 11580 12434 11608
rect 6932 11540 6960 11580
rect 6196 11512 6960 11540
rect 6089 11503 6147 11509
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7340 11512 7389 11540
rect 7340 11500 7346 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 9214 11540 9220 11552
rect 7800 11512 9220 11540
rect 7800 11500 7806 11512
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 11716 11549 11744 11580
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11509 11759 11543
rect 12406 11540 12434 11580
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 14200 11608 14228 11707
rect 12768 11580 14228 11608
rect 12768 11568 12774 11580
rect 14274 11540 14280 11552
rect 12406 11512 14280 11540
rect 11701 11503 11759 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14366 11500 14372 11552
rect 14424 11500 14430 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 1486 11336 1492 11348
rect 1443 11308 1492 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 2961 11339 3019 11345
rect 1596 11308 2176 11336
rect 1596 11141 1624 11308
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 1872 11064 1900 11231
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2038 11132 2044 11144
rect 1995 11104 2044 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2148 11132 2176 11308
rect 2961 11305 2973 11339
rect 3007 11336 3019 11339
rect 3142 11336 3148 11348
rect 3007 11308 3148 11336
rect 3007 11305 3019 11308
rect 2961 11299 3019 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 7374 11336 7380 11348
rect 4120 11308 7380 11336
rect 4120 11296 4126 11308
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7466 11296 7472 11348
rect 7524 11296 7530 11348
rect 8312 11308 8892 11336
rect 3602 11228 3608 11280
rect 3660 11268 3666 11280
rect 4157 11271 4215 11277
rect 4157 11268 4169 11271
rect 3660 11240 4169 11268
rect 3660 11228 3666 11240
rect 4157 11237 4169 11240
rect 4203 11237 4215 11271
rect 4157 11231 4215 11237
rect 5718 11228 5724 11280
rect 5776 11228 5782 11280
rect 6546 11228 6552 11280
rect 6604 11228 6610 11280
rect 7282 11228 7288 11280
rect 7340 11228 7346 11280
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 3237 11203 3295 11209
rect 2455 11172 3188 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2774 11132 2780 11144
rect 2148 11104 2780 11132
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 3160 11141 3188 11172
rect 3237 11169 3249 11203
rect 3283 11200 3295 11203
rect 3973 11203 4031 11209
rect 3973 11200 3985 11203
rect 3283 11172 3985 11200
rect 3283 11169 3295 11172
rect 3237 11163 3295 11169
rect 3973 11169 3985 11172
rect 4019 11169 4031 11203
rect 3973 11163 4031 11169
rect 3145 11135 3203 11141
rect 2832 11104 2912 11132
rect 2832 11092 2838 11104
rect 2884 11064 2912 11104
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 3191 11104 3617 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11132 3847 11135
rect 3835 11104 4016 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 1872 11036 2820 11064
rect 2884 11036 3188 11064
rect 2792 10996 2820 11036
rect 3160 11008 3188 11036
rect 3620 11008 3648 11095
rect 3988 11008 4016 11104
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4120 11104 4721 11132
rect 4120 11092 4126 11104
rect 4709 11101 4721 11104
rect 4755 11132 4767 11135
rect 5534 11132 5540 11144
rect 4755 11104 5540 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4798 11064 4804 11076
rect 4304 11036 4804 11064
rect 4304 11024 4310 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 4976 11067 5034 11073
rect 4976 11033 4988 11067
rect 5022 11064 5034 11067
rect 5736 11064 5764 11228
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6564 11200 6592 11228
rect 7300 11200 7328 11228
rect 6319 11172 6592 11200
rect 6932 11172 7328 11200
rect 7484 11200 7512 11296
rect 7653 11271 7711 11277
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7742 11268 7748 11280
rect 7699 11240 7748 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7837 11271 7895 11277
rect 7837 11237 7849 11271
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 8113 11271 8171 11277
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 8312 11268 8340 11308
rect 8159 11240 8340 11268
rect 8864 11268 8892 11308
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8996 11308 9321 11336
rect 8996 11296 9002 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 9309 11299 9367 11305
rect 9646 11308 11468 11336
rect 8864 11240 9168 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 7852 11200 7880 11231
rect 9140 11209 9168 11240
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 9646 11268 9674 11308
rect 9272 11240 9674 11268
rect 11440 11268 11468 11308
rect 11882 11296 11888 11348
rect 11940 11296 11946 11348
rect 13262 11336 13268 11348
rect 12406 11308 13268 11336
rect 12406 11268 12434 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13630 11296 13636 11348
rect 13688 11296 13694 11348
rect 11440 11240 12434 11268
rect 9272 11228 9278 11240
rect 9125 11203 9183 11209
rect 7484 11172 7788 11200
rect 7852 11172 8340 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6932 11132 6960 11172
rect 6503 11104 6960 11132
rect 7760 11132 7788 11172
rect 8312 11141 8340 11172
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11940 11172 11989 11200
rect 11940 11160 11946 11172
rect 11977 11169 11989 11172
rect 12023 11200 12035 11203
rect 13081 11203 13139 11209
rect 12023 11172 12434 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7760 11104 8033 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 5022 11036 5764 11064
rect 5022 11033 5034 11036
rect 4976 11027 5034 11033
rect 6822 11024 6828 11076
rect 6880 11024 6886 11076
rect 6917 11067 6975 11073
rect 6917 11033 6929 11067
rect 6963 11064 6975 11067
rect 7098 11064 7104 11076
rect 6963 11036 7104 11064
rect 6963 11033 6975 11036
rect 6917 11027 6975 11033
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7193 11067 7251 11073
rect 7193 11033 7205 11067
rect 7239 11033 7251 11067
rect 8036 11064 8064 11095
rect 8404 11064 8432 11095
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8904 11104 8953 11132
rect 8904 11092 8910 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11132 10563 11135
rect 11054 11132 11060 11144
rect 10551 11104 11060 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12406 11132 12434 11172
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 13648 11200 13676 11296
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13780 11240 14105 11268
rect 13780 11228 13786 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 13127 11172 13676 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12406 11104 12725 11132
rect 12713 11101 12725 11104
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 14274 11092 14280 11144
rect 14332 11092 14338 11144
rect 8036 11036 8432 11064
rect 8496 11064 8524 11092
rect 10410 11064 10416 11076
rect 8496 11036 10416 11064
rect 7193 11027 7251 11033
rect 3050 10996 3056 11008
rect 2792 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 3142 10956 3148 11008
rect 3200 10956 3206 11008
rect 3602 10956 3608 11008
rect 3660 10956 3666 11008
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 5592 10968 6101 10996
rect 5592 10956 5598 10968
rect 6089 10965 6101 10968
rect 6135 10965 6147 10999
rect 6840 10996 6868 11024
rect 7208 10996 7236 11027
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 10772 11067 10830 11073
rect 10772 11033 10784 11067
rect 10818 11064 10830 11067
rect 12176 11064 12204 11092
rect 10818 11036 12204 11064
rect 13173 11067 13231 11073
rect 10818 11033 10830 11036
rect 10772 11027 10830 11033
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13354 11064 13360 11076
rect 13219 11036 13360 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 13648 11036 13737 11064
rect 13648 11008 13676 11036
rect 13725 11033 13737 11036
rect 13771 11033 13783 11067
rect 13725 11027 13783 11033
rect 6840 10968 7236 10996
rect 6089 10959 6147 10965
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10686 10996 10692 11008
rect 10008 10968 10692 10996
rect 10008 10956 10014 10968
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 12802 10956 12808 11008
rect 12860 10956 12866 11008
rect 13630 10956 13636 11008
rect 13688 10956 13694 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3326 10792 3332 10804
rect 2915 10764 3332 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 4062 10752 4068 10804
rect 4120 10752 4126 10804
rect 5166 10752 5172 10804
rect 5224 10752 5230 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5994 10792 6000 10804
rect 5307 10764 6000 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7837 10795 7895 10801
rect 7837 10792 7849 10795
rect 7156 10764 7849 10792
rect 7156 10752 7162 10764
rect 7837 10761 7849 10764
rect 7883 10761 7895 10795
rect 7837 10755 7895 10761
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 8846 10792 8852 10804
rect 8527 10764 8852 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8996 10764 9321 10792
rect 8996 10752 9002 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 12158 10792 12164 10804
rect 9456 10764 12164 10792
rect 9456 10752 9462 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13495 10764 13952 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 4080 10724 4108 10752
rect 6181 10727 6239 10733
rect 6181 10724 6193 10727
rect 3804 10696 4108 10724
rect 5092 10696 6193 10724
rect 3804 10668 3832 10696
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 992 10628 1593 10656
rect 992 10616 998 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 1946 10616 1952 10668
rect 2004 10616 2010 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1728 10560 2145 10588
rect 1728 10548 1734 10560
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10557 2375 10591
rect 3068 10588 3096 10619
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3292 10628 3617 10656
rect 3292 10616 3298 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 4056 10659 4114 10665
rect 4056 10625 4068 10659
rect 4102 10656 4114 10659
rect 5092 10656 5120 10696
rect 6181 10693 6193 10696
rect 6227 10693 6239 10727
rect 6181 10687 6239 10693
rect 6546 10684 6552 10736
rect 6604 10684 6610 10736
rect 7650 10684 7656 10736
rect 7708 10684 7714 10736
rect 8754 10724 8760 10736
rect 8404 10696 8760 10724
rect 4102 10628 5120 10656
rect 5445 10659 5503 10665
rect 4102 10625 4114 10628
rect 4056 10619 4114 10625
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7668 10656 7696 10684
rect 8404 10665 8432 10696
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 8864 10724 8892 10752
rect 11876 10727 11934 10733
rect 8864 10696 9444 10724
rect 7147 10628 7696 10656
rect 7929 10659 7987 10665
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 3326 10588 3332 10600
rect 3068 10560 3332 10588
rect 2317 10551 2375 10557
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 2332 10520 2360 10551
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 1811 10492 2360 10520
rect 2777 10523 2835 10529
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 2777 10489 2789 10523
rect 2823 10520 2835 10523
rect 5460 10520 5488 10619
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 6454 10588 6460 10600
rect 5629 10551 5687 10557
rect 6012 10560 6460 10588
rect 2823 10492 3740 10520
rect 5460 10492 5580 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 1394 10412 1400 10464
rect 1452 10412 1458 10464
rect 3234 10412 3240 10464
rect 3292 10412 3298 10464
rect 3418 10412 3424 10464
rect 3476 10412 3482 10464
rect 3712 10452 3740 10492
rect 5552 10464 5580 10492
rect 3970 10452 3976 10464
rect 3712 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 5644 10452 5672 10551
rect 6012 10532 6040 10560
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7340 10560 7389 10588
rect 7340 10548 7346 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 5994 10480 6000 10532
rect 6052 10480 6058 10532
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7944 10520 7972 10619
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 9416 10665 9444 10696
rect 9508 10696 11744 10724
rect 8849 10659 8907 10665
rect 8849 10656 8861 10659
rect 8536 10628 8861 10656
rect 8536 10616 8542 10628
rect 8849 10625 8861 10628
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9214 10588 9220 10600
rect 8711 10560 9220 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 7156 10492 7972 10520
rect 8113 10523 8171 10529
rect 7156 10480 7162 10492
rect 8113 10489 8125 10523
rect 8159 10520 8171 10523
rect 9508 10520 9536 10696
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 10100 10628 10149 10656
rect 10100 10616 10106 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10560 10628 10609 10656
rect 10560 10616 10566 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 10643 10628 11008 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9585 10551 9643 10557
rect 9968 10560 10241 10588
rect 8159 10492 9536 10520
rect 8159 10489 8171 10492
rect 8113 10483 8171 10489
rect 6730 10452 6736 10464
rect 5644 10424 6736 10452
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9600 10452 9628 10551
rect 9968 10464 9996 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 10275 10560 10701 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10689 10557 10701 10560
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 10980 10588 11008 10628
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11606 10656 11612 10668
rect 11112 10628 11612 10656
rect 11112 10616 11118 10628
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 11716 10656 11744 10696
rect 11876 10693 11888 10727
rect 11922 10724 11934 10727
rect 12618 10724 12624 10736
rect 11922 10696 12624 10724
rect 11922 10693 11934 10696
rect 11876 10687 11934 10693
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 13924 10733 13952 10764
rect 13909 10727 13967 10733
rect 13228 10696 13400 10724
rect 13228 10684 13234 10696
rect 13372 10656 13400 10696
rect 13909 10693 13921 10727
rect 13955 10693 13967 10727
rect 13909 10687 13967 10693
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 11716 10628 13308 10656
rect 13372 10628 13645 10656
rect 11146 10588 11152 10600
rect 10980 10560 11152 10588
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 13280 10520 13308 10628
rect 13633 10625 13645 10628
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13504 10560 13829 10588
rect 13504 10548 13510 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 13280 10492 13584 10520
rect 9456 10424 9628 10452
rect 9456 10412 9462 10424
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 10410 10412 10416 10464
rect 10468 10412 10474 10464
rect 11330 10412 11336 10464
rect 11388 10412 11394 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12768 10424 13001 10452
rect 12768 10412 12774 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 13556 10452 13584 10492
rect 13630 10480 13636 10532
rect 13688 10520 13694 10532
rect 14108 10520 14136 10551
rect 13688 10492 14136 10520
rect 13688 10480 13694 10492
rect 14090 10452 14096 10464
rect 13556 10424 14096 10452
rect 12989 10415 13047 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 3786 10248 3792 10260
rect 1504 10220 3792 10248
rect 1504 10121 1532 10220
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4028 10220 4169 10248
rect 4028 10208 4034 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5994 10248 6000 10260
rect 5215 10220 6000 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6178 10208 6184 10260
rect 6236 10248 6242 10260
rect 6236 10220 6500 10248
rect 6236 10208 6242 10220
rect 3418 10140 3424 10192
rect 3476 10180 3482 10192
rect 4890 10180 4896 10192
rect 3476 10152 4896 10180
rect 3476 10140 3482 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 6362 10180 6368 10192
rect 5920 10152 6368 10180
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10081 1547 10115
rect 1489 10075 1547 10081
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3191 10084 3985 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5920 10112 5948 10152
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 4755 10084 5948 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5994 10072 6000 10124
rect 6052 10072 6058 10124
rect 6086 10072 6092 10124
rect 6144 10112 6150 10124
rect 6472 10112 6500 10220
rect 6546 10208 6552 10260
rect 6604 10208 6610 10260
rect 6825 10251 6883 10257
rect 6825 10217 6837 10251
rect 6871 10248 6883 10251
rect 7282 10248 7288 10260
rect 6871 10220 7288 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 9646 10220 9904 10248
rect 6564 10180 6592 10208
rect 7101 10183 7159 10189
rect 7101 10180 7113 10183
rect 6564 10152 7113 10180
rect 7101 10149 7113 10152
rect 7147 10149 7159 10183
rect 9416 10180 9444 10208
rect 9493 10183 9551 10189
rect 9493 10180 9505 10183
rect 9416 10152 9505 10180
rect 7101 10143 7159 10149
rect 9493 10149 9505 10152
rect 9539 10149 9551 10183
rect 9493 10143 9551 10149
rect 6914 10112 6920 10124
rect 6144 10084 6316 10112
rect 6472 10084 6920 10112
rect 6144 10072 6150 10084
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3694 10044 3700 10056
rect 3375 10016 3700 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 3878 10044 3884 10056
rect 3835 10016 3884 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4304 10016 4537 10044
rect 4304 10004 4310 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 1756 9979 1814 9985
rect 1756 9945 1768 9979
rect 1802 9976 1814 9979
rect 2130 9976 2136 9988
rect 1802 9948 2136 9976
rect 1802 9945 1814 9948
rect 1756 9939 1814 9945
rect 2130 9936 2136 9948
rect 2188 9936 2194 9988
rect 5368 9976 5396 10007
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5776 10016 6193 10044
rect 5776 10004 5782 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6288 10044 6316 10084
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 9214 10072 9220 10124
rect 9272 10112 9278 10124
rect 9646 10112 9674 10220
rect 9876 10180 9904 10220
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 10100 10220 10149 10248
rect 10100 10208 10106 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10870 10248 10876 10260
rect 10551 10220 10876 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 11388 10220 11897 10248
rect 11388 10208 11394 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 11885 10211 11943 10217
rect 9876 10152 10088 10180
rect 9272 10084 9674 10112
rect 9272 10072 9278 10084
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 10060 10112 10088 10152
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 10652 10152 11437 10180
rect 10652 10140 10658 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 10060 10084 10364 10112
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6288 10016 6745 10044
rect 6181 10007 6239 10013
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 5534 9976 5540 9988
rect 2884 9948 3648 9976
rect 5368 9948 5540 9976
rect 2884 9917 2912 9948
rect 3620 9920 3648 9948
rect 5534 9936 5540 9948
rect 5592 9976 5598 9988
rect 7024 9976 7052 10007
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9306 10044 9312 10056
rect 9171 10016 9312 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9674 10044 9680 10056
rect 9447 10016 9680 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9876 10016 9965 10044
rect 5592 9948 7052 9976
rect 7552 9979 7610 9985
rect 5592 9936 5598 9948
rect 7552 9945 7564 9979
rect 7598 9976 7610 9979
rect 9766 9976 9772 9988
rect 7598 9948 9772 9976
rect 7598 9945 7610 9948
rect 7552 9939 7610 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9877 2927 9911
rect 2869 9871 2927 9877
rect 3418 9868 3424 9920
rect 3476 9868 3482 9920
rect 3602 9868 3608 9920
rect 3660 9868 3666 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5408 9880 5917 9908
rect 5408 9868 5414 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6052 9880 6653 9908
rect 6052 9868 6058 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 6641 9871 6699 9877
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 6788 9880 8677 9908
rect 6788 9868 6794 9880
rect 8665 9877 8677 9880
rect 8711 9877 8723 9911
rect 8665 9871 8723 9877
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9876 9908 9904 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 9456 9880 9904 9908
rect 10336 9908 10364 10084
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11517 10115 11575 10121
rect 10468 10084 10732 10112
rect 10468 10072 10474 10084
rect 10704 10053 10732 10084
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11900 10112 11928 10211
rect 14366 10208 14372 10260
rect 14424 10208 14430 10260
rect 12897 10183 12955 10189
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 13446 10180 13452 10192
rect 12943 10152 13452 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11563 10084 11836 10112
rect 11900 10084 12265 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 10888 9976 10916 10007
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11808 10044 11836 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 12802 10112 12808 10124
rect 12483 10084 12808 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13722 10112 13728 10124
rect 13311 10084 13728 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 11974 10044 11980 10056
rect 11808 10016 11980 10044
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 12216 10016 13032 10044
rect 12216 10004 12222 10016
rect 12710 9976 12716 9988
rect 10888 9948 12716 9976
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 12894 9936 12900 9988
rect 12952 9936 12958 9988
rect 13004 9976 13032 10016
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13228 10016 14197 10044
rect 13228 10004 13234 10016
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 14476 9976 14504 10004
rect 13004 9948 14504 9976
rect 10962 9908 10968 9920
rect 10336 9880 10968 9908
rect 9456 9868 9462 9880
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12618 9908 12624 9920
rect 12216 9880 12624 9908
rect 12216 9868 12222 9880
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12912 9908 12940 9936
rect 13630 9908 13636 9920
rect 12912 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 1394 9664 1400 9716
rect 1452 9664 1458 9716
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9704 1639 9707
rect 1670 9704 1676 9716
rect 1627 9676 1676 9704
rect 1627 9673 1639 9676
rect 1581 9667 1639 9673
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 1765 9707 1823 9713
rect 1765 9673 1777 9707
rect 1811 9704 1823 9707
rect 1946 9704 1952 9716
rect 1811 9676 1952 9704
rect 1811 9673 1823 9676
rect 1765 9667 1823 9673
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 3694 9704 3700 9716
rect 3200 9676 3700 9704
rect 3200 9664 3206 9676
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 3878 9664 3884 9716
rect 3936 9664 3942 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4304 9676 4629 9704
rect 4304 9664 4310 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4617 9667 4675 9673
rect 5166 9664 5172 9716
rect 5224 9664 5230 9716
rect 5997 9707 6055 9713
rect 5997 9673 6009 9707
rect 6043 9704 6055 9707
rect 6178 9704 6184 9716
rect 6043 9676 6184 9704
rect 6043 9673 6055 9676
rect 5997 9667 6055 9673
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6454 9704 6460 9716
rect 6380 9676 6460 9704
rect 6380 9674 6408 9676
rect 1412 9568 1440 9664
rect 3896 9636 3924 9664
rect 5184 9636 5212 9664
rect 6288 9646 6408 9674
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 7469 9707 7527 9713
rect 6604 9676 6960 9704
rect 6604 9664 6610 9676
rect 5905 9639 5963 9645
rect 1964 9608 3096 9636
rect 3896 9608 4016 9636
rect 1964 9577 1992 9608
rect 3068 9580 3096 9608
rect 1489 9571 1547 9577
rect 1489 9568 1501 9571
rect 1412 9540 1501 9568
rect 1489 9537 1501 9540
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2406 9528 2412 9580
rect 2464 9528 2470 9580
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3988 9577 4016 9608
rect 5000 9608 5580 9636
rect 5000 9577 5028 9608
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3476 9540 3617 9568
rect 3476 9528 3482 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4939 9540 4997 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5123 9540 5457 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5552 9568 5580 9608
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 6288 9636 6316 9646
rect 5951 9608 6316 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 6730 9596 6736 9648
rect 6788 9596 6794 9648
rect 6932 9636 6960 9676
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7515 9676 7549 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 6932 9608 7043 9636
rect 5994 9568 6000 9580
rect 5552 9540 6000 9568
rect 5445 9531 5503 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 2501 9503 2559 9509
rect 2501 9500 2513 9503
rect 1728 9472 2513 9500
rect 1728 9460 1734 9472
rect 2501 9469 2513 9472
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9469 2743 9503
rect 3142 9500 3148 9512
rect 2685 9463 2743 9469
rect 3068 9472 3148 9500
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2700 9432 2728 9463
rect 2271 9404 2728 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 3068 9364 3096 9472
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3896 9500 3924 9531
rect 5994 9528 6000 9540
rect 6052 9558 6058 9580
rect 6189 9571 6247 9577
rect 6189 9558 6201 9571
rect 6052 9537 6201 9558
rect 6235 9537 6247 9571
rect 6052 9531 6247 9537
rect 6052 9530 6224 9531
rect 6052 9528 6058 9530
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6748 9568 6776 9596
rect 6687 9540 6776 9568
rect 6917 9571 6975 9577
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 3436 9472 3924 9500
rect 4157 9503 4215 9509
rect 3436 9441 3464 9472
rect 4157 9469 4169 9503
rect 4203 9469 4215 9503
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 4157 9463 4215 9469
rect 4632 9472 5273 9500
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9401 3479 9435
rect 3421 9395 3479 9401
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4172 9432 4200 9463
rect 3743 9404 4200 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 1820 9336 3096 9364
rect 3145 9367 3203 9373
rect 1820 9324 1826 9336
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 4632 9364 4660 9472
rect 5261 9469 5273 9472
rect 5307 9500 5319 9503
rect 5902 9500 5908 9512
rect 5307 9472 5908 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6380 9441 6408 9528
rect 6564 9500 6592 9531
rect 6472 9472 6592 9500
rect 4709 9435 4767 9441
rect 4709 9401 4721 9435
rect 4755 9432 4767 9435
rect 6365 9435 6423 9441
rect 4755 9404 6224 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 3191 9336 4660 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5902 9364 5908 9376
rect 5132 9336 5908 9364
rect 5132 9324 5138 9336
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6196 9364 6224 9404
rect 6365 9401 6377 9435
rect 6411 9401 6423 9435
rect 6365 9395 6423 9401
rect 6472 9364 6500 9472
rect 6196 9336 6500 9364
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6656 9364 6684 9531
rect 6730 9460 6736 9512
rect 6788 9460 6794 9512
rect 6748 9432 6776 9460
rect 6932 9444 6960 9531
rect 6748 9404 6868 9432
rect 6604 9336 6684 9364
rect 6604 9324 6610 9336
rect 6730 9324 6736 9376
rect 6788 9324 6794 9376
rect 6840 9364 6868 9404
rect 6914 9392 6920 9444
rect 6972 9392 6978 9444
rect 7015 9432 7043 9608
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7285 9639 7343 9645
rect 7285 9636 7297 9639
rect 7156 9608 7297 9636
rect 7156 9596 7162 9608
rect 7285 9605 7297 9608
rect 7331 9605 7343 9639
rect 7484 9636 7512 9667
rect 9398 9664 9404 9716
rect 9456 9704 9462 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 9456 9676 9781 9704
rect 9456 9664 9462 9676
rect 9769 9673 9781 9676
rect 9815 9673 9827 9707
rect 9769 9667 9827 9673
rect 11698 9664 11704 9716
rect 11756 9664 11762 9716
rect 12158 9664 12164 9716
rect 12216 9664 12222 9716
rect 12894 9704 12900 9716
rect 12636 9676 12900 9704
rect 9030 9636 9036 9648
rect 7484 9608 9036 9636
rect 7285 9599 7343 9605
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 12636 9636 12664 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 12989 9707 13047 9713
rect 12989 9673 13001 9707
rect 13035 9704 13047 9707
rect 13078 9704 13084 9716
rect 13035 9676 13084 9704
rect 13035 9673 13047 9676
rect 12989 9667 13047 9673
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 14182 9664 14188 9716
rect 14240 9664 14246 9716
rect 10560 9608 11100 9636
rect 10560 9596 10566 9608
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 7101 9435 7159 9441
rect 7101 9432 7113 9435
rect 7015 9404 7113 9432
rect 7101 9401 7113 9404
rect 7147 9401 7159 9435
rect 7101 9395 7159 9401
rect 7208 9364 7236 9531
rect 7668 9444 7696 9531
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9669 9571 9727 9577
rect 8895 9540 9628 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8294 9500 8300 9512
rect 8251 9472 8300 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8496 9500 8524 9531
rect 9122 9500 9128 9512
rect 8496 9472 9128 9500
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 7650 9392 7656 9444
rect 7708 9392 7714 9444
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9306 9432 9312 9444
rect 8628 9404 9312 9432
rect 8628 9392 8634 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9490 9392 9496 9444
rect 9548 9392 9554 9444
rect 6840 9336 7236 9364
rect 7926 9324 7932 9376
rect 7984 9324 7990 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 8720 9336 9413 9364
rect 8720 9324 8726 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9600 9364 9628 9540
rect 9669 9537 9681 9571
rect 9715 9568 9727 9571
rect 9766 9568 9772 9580
rect 9715 9540 9772 9568
rect 9715 9537 9727 9540
rect 9669 9531 9727 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9876 9540 9965 9568
rect 9876 9500 9904 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10183 9540 10272 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 9784 9472 9904 9500
rect 9784 9444 9812 9472
rect 9766 9392 9772 9444
rect 9824 9392 9830 9444
rect 10060 9376 10088 9531
rect 10042 9364 10048 9376
rect 9600 9336 10048 9364
rect 9401 9327 9459 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10244 9364 10272 9540
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10468 9540 10793 9568
rect 10468 9528 10474 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 10318 9460 10324 9512
rect 10376 9460 10382 9512
rect 11072 9500 11100 9608
rect 11164 9608 12664 9636
rect 11164 9577 11192 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 12768 9608 13308 9636
rect 12768 9596 12774 9608
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11296 9540 11621 9568
rect 11296 9528 11302 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 12345 9571 12403 9577
rect 12345 9558 12357 9571
rect 11885 9531 11943 9537
rect 12259 9537 12357 9558
rect 12391 9537 12403 9571
rect 12259 9531 12403 9537
rect 11698 9500 11704 9512
rect 11072 9472 11704 9500
rect 11698 9460 11704 9472
rect 11756 9500 11762 9512
rect 11900 9500 11928 9531
rect 12259 9530 12388 9531
rect 11756 9472 11928 9500
rect 11756 9460 11762 9472
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12259 9500 12287 9530
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13280 9577 13308 9608
rect 13354 9596 13360 9648
rect 13412 9596 13418 9648
rect 13464 9608 14412 9636
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12860 9540 12909 9568
rect 12860 9528 12866 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13464 9568 13492 9608
rect 13311 9540 13492 9568
rect 13725 9571 13783 9577
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13740 9500 13768 9531
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 14384 9577 14412 9608
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 12216 9472 12287 9500
rect 12452 9472 13768 9500
rect 12216 9460 12222 9472
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 12452 9441 12480 9472
rect 10597 9435 10655 9441
rect 10597 9432 10609 9435
rect 10468 9404 10609 9432
rect 10468 9392 10474 9404
rect 10597 9401 10609 9404
rect 10643 9401 10655 9435
rect 12437 9435 12495 9441
rect 10597 9395 10655 9401
rect 10980 9404 12296 9432
rect 10502 9364 10508 9376
rect 10244 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10980 9373 11008 9404
rect 10965 9367 11023 9373
rect 10965 9333 10977 9367
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 11241 9367 11299 9373
rect 11241 9333 11253 9367
rect 11287 9364 11299 9367
rect 11882 9364 11888 9376
rect 11287 9336 11888 9364
rect 11287 9333 11299 9336
rect 11241 9327 11299 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11974 9324 11980 9376
rect 12032 9324 12038 9376
rect 12268 9364 12296 9404
rect 12437 9401 12449 9435
rect 12483 9401 12495 9435
rect 12437 9395 12495 9401
rect 12636 9404 13860 9432
rect 12636 9364 12664 9404
rect 13832 9376 13860 9404
rect 12268 9336 12664 9364
rect 12713 9367 12771 9373
rect 12713 9333 12725 9367
rect 12759 9364 12771 9367
rect 13354 9364 13360 9376
rect 12759 9336 13360 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13814 9324 13820 9376
rect 13872 9324 13878 9376
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 2406 9160 2412 9172
rect 2179 9132 2412 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3053 9163 3111 9169
rect 3053 9160 3065 9163
rect 2740 9132 3065 9160
rect 2740 9120 2746 9132
rect 3053 9129 3065 9132
rect 3099 9129 3111 9163
rect 3053 9123 3111 9129
rect 3142 9120 3148 9172
rect 3200 9160 3206 9172
rect 3970 9160 3976 9172
rect 3200 9132 3976 9160
rect 3200 9120 3206 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 4246 9120 4252 9172
rect 4304 9120 4310 9172
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5031 9132 5672 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 3418 9052 3424 9104
rect 3476 9052 3482 9104
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9061 5319 9095
rect 5644 9092 5672 9132
rect 5718 9120 5724 9172
rect 5776 9120 5782 9172
rect 6012 9132 6960 9160
rect 6012 9104 6040 9132
rect 5994 9092 6000 9104
rect 5644 9064 6000 9092
rect 5261 9055 5319 9061
rect 3436 9024 3464 9052
rect 2332 8996 3464 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 992 8928 1593 8956
rect 992 8916 998 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 1872 8888 1900 8919
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 2332 8965 2360 8996
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 3436 8965 3464 8996
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3559 8996 3985 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 5276 9024 5304 9055
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 6932 9092 6960 9132
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7650 9160 7656 9172
rect 7300 9132 7656 9160
rect 7300 9092 7328 9132
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8352 9132 10548 9160
rect 8352 9120 8358 9132
rect 6135 9064 6868 9092
rect 6932 9064 7328 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 6457 9027 6515 9033
rect 5276 8996 6408 9024
rect 3973 8987 4031 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2870 8959 2928 8965
rect 2870 8925 2882 8959
rect 2916 8925 2928 8959
rect 2870 8919 2928 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 952 8860 1900 8888
rect 2240 8888 2268 8916
rect 2700 8888 2728 8919
rect 2240 8860 2728 8888
rect 2884 8888 2912 8919
rect 3142 8888 3148 8900
rect 2884 8860 3148 8888
rect 952 8832 980 8860
rect 934 8780 940 8832
rect 992 8780 998 8832
rect 1394 8780 1400 8832
rect 1452 8780 1458 8832
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8820 2099 8823
rect 2314 8820 2320 8832
rect 2087 8792 2320 8820
rect 2087 8789 2099 8792
rect 2041 8783 2099 8789
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 2406 8780 2412 8832
rect 2464 8780 2470 8832
rect 2700 8820 2728 8860
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3804 8820 3832 8919
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4816 8888 4844 8919
rect 5074 8916 5080 8968
rect 5132 8916 5138 8968
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8932 5411 8959
rect 5399 8925 5488 8932
rect 5353 8919 5488 8925
rect 5376 8904 5488 8919
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6380 8965 6408 8996
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6638 9024 6644 9036
rect 6503 8996 6644 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 6840 9033 6868 9064
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 10100 9064 10333 9092
rect 10100 9052 10106 9064
rect 10321 9061 10333 9064
rect 10367 9061 10379 9095
rect 10520 9092 10548 9132
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12618 9160 12624 9172
rect 11756 9132 12624 9160
rect 11756 9120 11762 9132
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 10520 9064 10640 9092
rect 10321 9055 10379 9061
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 10612 9024 10640 9064
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 14090 9092 14096 9104
rect 11020 9064 12020 9092
rect 11020 9052 11026 9064
rect 11146 9024 11152 9036
rect 10612 8996 11152 9024
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11992 9033 12020 9064
rect 12406 9064 14096 9092
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 9024 12219 9027
rect 12406 9024 12434 9064
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 14366 9052 14372 9104
rect 14424 9052 14430 9104
rect 12207 8996 12434 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 13354 8984 13360 9036
rect 13412 8984 13418 9036
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8956 6423 8959
rect 6411 8928 6868 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 5166 8888 5172 8900
rect 4816 8860 5172 8888
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 5460 8888 5488 8904
rect 5644 8888 5672 8916
rect 6840 8900 6868 8928
rect 6546 8888 6552 8900
rect 5460 8860 5580 8888
rect 5644 8860 6552 8888
rect 2700 8792 3832 8820
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4304 8792 4537 8820
rect 4304 8780 4310 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 5552 8820 5580 8860
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 6822 8848 6828 8900
rect 6880 8848 6886 8900
rect 6362 8820 6368 8832
rect 5552 8792 6368 8820
rect 6362 8780 6368 8792
rect 6420 8820 6426 8832
rect 6932 8820 6960 8984
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 7340 8928 7389 8956
rect 7340 8916 7346 8928
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 7423 8928 8953 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 11241 8959 11299 8965
rect 8987 8928 9444 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9416 8900 9444 8928
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 7644 8891 7702 8897
rect 7644 8857 7656 8891
rect 7690 8888 7702 8891
rect 8662 8888 8668 8900
rect 7690 8860 8668 8888
rect 7690 8857 7702 8860
rect 7644 8851 7702 8857
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 9208 8891 9266 8897
rect 9208 8857 9220 8891
rect 9254 8888 9266 8891
rect 9254 8860 9352 8888
rect 9254 8857 9266 8860
rect 9208 8851 9266 8857
rect 6420 8792 6960 8820
rect 6420 8780 6426 8792
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8757 8823 8815 8829
rect 8757 8820 8769 8823
rect 7800 8792 8769 8820
rect 7800 8780 7806 8792
rect 8757 8789 8769 8792
rect 8803 8789 8815 8823
rect 9324 8820 9352 8860
rect 9398 8848 9404 8900
rect 9456 8848 9462 8900
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 11149 8891 11207 8897
rect 11149 8888 11161 8891
rect 10980 8860 11161 8888
rect 9766 8820 9772 8832
rect 9324 8792 9772 8820
rect 8757 8783 8815 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10980 8820 11008 8860
rect 11149 8857 11161 8860
rect 11195 8857 11207 8891
rect 11149 8851 11207 8857
rect 10560 8792 11008 8820
rect 10560 8780 10566 8792
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11256 8820 11284 8919
rect 11882 8916 11888 8968
rect 11940 8916 11946 8968
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8956 12863 8959
rect 12894 8956 12900 8968
rect 12851 8928 12900 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13372 8956 13400 8984
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 13372 8928 13645 8956
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 13722 8916 13728 8968
rect 13780 8916 13786 8968
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8925 14243 8959
rect 14185 8919 14243 8925
rect 11900 8888 11928 8916
rect 14200 8888 14228 8919
rect 11900 8860 14228 8888
rect 11112 8792 11284 8820
rect 11112 8780 11118 8792
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 12618 8780 12624 8832
rect 12676 8780 12682 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 12860 8792 13369 8820
rect 12860 8780 12866 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 13357 8783 13415 8789
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13596 8792 13921 8820
rect 13596 8780 13602 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 2188 8588 3433 8616
rect 2188 8576 2194 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 4982 8616 4988 8628
rect 4724 8588 4988 8616
rect 3602 8548 3608 8560
rect 2516 8520 3608 8548
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 2516 8424 2544 8520
rect 3602 8508 3608 8520
rect 3660 8548 3666 8560
rect 3660 8520 4292 8548
rect 3660 8508 3666 8520
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2682 8480 2688 8492
rect 2639 8452 2688 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2682 8440 2688 8452
rect 2740 8484 2746 8492
rect 2740 8480 2774 8484
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 2740 8452 3525 8480
rect 2740 8440 2746 8452
rect 3513 8449 3525 8452
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 4264 8489 4292 8520
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 4724 8480 4752 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 6328 8588 6377 8616
rect 6328 8576 6334 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 7248 8588 7297 8616
rect 7248 8576 7254 8588
rect 7285 8585 7297 8588
rect 7331 8585 7343 8619
rect 7285 8579 7343 8585
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9950 8616 9956 8628
rect 9723 8588 9956 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10318 8616 10324 8628
rect 10060 8588 10324 8616
rect 4792 8551 4850 8557
rect 4792 8517 4804 8551
rect 4838 8548 4850 8551
rect 5350 8548 5356 8560
rect 4838 8520 5356 8548
rect 4838 8517 4850 8520
rect 4792 8511 4850 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 6454 8508 6460 8560
rect 6512 8548 6518 8560
rect 6748 8548 6776 8576
rect 6512 8520 6684 8548
rect 6748 8520 6868 8548
rect 6512 8508 6518 8520
rect 4672 8452 5580 8480
rect 4672 8440 4678 8452
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1728 8384 1961 8412
rect 1728 8372 1734 8384
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 2130 8372 2136 8424
rect 2188 8372 2194 8424
rect 2498 8372 2504 8424
rect 2556 8372 2562 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3050 8412 3056 8424
rect 2915 8384 3056 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 3804 8412 3832 8440
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 3804 8384 4537 8412
rect 3697 8375 3755 8381
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 1762 8344 1768 8356
rect 1627 8316 1768 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 3712 8344 3740 8375
rect 3878 8344 3884 8356
rect 3712 8316 3884 8344
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 5552 8344 5580 8452
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6656 8480 6684 8520
rect 6730 8480 6736 8492
rect 6656 8452 6736 8480
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6840 8489 6868 8520
rect 7374 8508 7380 8560
rect 7432 8508 7438 8560
rect 10060 8557 10088 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10410 8576 10416 8628
rect 10468 8576 10474 8628
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10836 8588 10885 8616
rect 10836 8576 10842 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 12618 8576 12624 8628
rect 12676 8576 12682 8628
rect 12894 8576 12900 8628
rect 12952 8576 12958 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 13096 8588 14473 8616
rect 10045 8551 10103 8557
rect 7484 8520 9674 8548
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 7484 8480 7512 8520
rect 9646 8492 9674 8520
rect 10045 8517 10057 8551
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 10428 8548 10456 8576
rect 10183 8520 10456 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 11716 8548 11744 8576
rect 10560 8520 11744 8548
rect 11784 8551 11842 8557
rect 10560 8508 10566 8520
rect 11784 8517 11796 8551
rect 11830 8548 11842 8551
rect 11900 8548 11928 8576
rect 11830 8520 11928 8548
rect 12636 8548 12664 8576
rect 13096 8557 13124 8588
rect 14461 8585 14473 8588
rect 14507 8585 14519 8619
rect 14461 8579 14519 8585
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 12636 8520 13093 8548
rect 11830 8517 11842 8520
rect 11784 8511 11842 8517
rect 13081 8517 13093 8520
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 13173 8551 13231 8557
rect 13173 8517 13185 8551
rect 13219 8548 13231 8551
rect 14366 8548 14372 8560
rect 13219 8520 14372 8548
rect 13219 8517 13231 8520
rect 13173 8511 13231 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 6825 8443 6883 8449
rect 6932 8452 7512 8480
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6512 8384 6653 8412
rect 6512 8372 6518 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 6932 8344 6960 8452
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 8352 8452 9413 8480
rect 8352 8440 8358 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9646 8452 9680 8492
rect 9401 8443 9459 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10836 8452 11069 8480
rect 10836 8440 10842 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11606 8480 11612 8492
rect 11563 8452 11612 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 11164 8412 11192 8443
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 12894 8440 12900 8492
rect 12952 8440 12958 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 7064 8400 10732 8412
rect 10888 8400 11192 8412
rect 7064 8384 11192 8400
rect 12912 8412 12940 8440
rect 13906 8412 13912 8424
rect 12912 8384 13912 8412
rect 7064 8372 7070 8384
rect 10704 8372 10916 8384
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14182 8412 14188 8424
rect 14047 8384 14188 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 4028 8316 4568 8344
rect 5552 8316 6960 8344
rect 7015 8316 8800 8344
rect 4028 8304 4034 8316
rect 4338 8236 4344 8288
rect 4396 8236 4402 8288
rect 4540 8276 4568 8316
rect 5626 8276 5632 8288
rect 4540 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 7015 8276 7043 8316
rect 8772 8288 8800 8316
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 10502 8344 10508 8356
rect 8996 8316 10508 8344
rect 8996 8304 9002 8316
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 10594 8304 10600 8356
rect 10652 8304 10658 8356
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11204 8316 11468 8344
rect 11204 8304 11210 8316
rect 5960 8248 7043 8276
rect 5960 8236 5966 8248
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8260 8248 8677 8276
rect 8260 8236 8266 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 8754 8236 8760 8288
rect 8812 8236 8818 8288
rect 9214 8236 9220 8288
rect 9272 8236 9278 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 10778 8276 10784 8288
rect 9732 8248 10784 8276
rect 9732 8236 9738 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11330 8236 11336 8288
rect 11388 8236 11394 8288
rect 11440 8276 11468 8316
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 13596 8316 13645 8344
rect 13596 8304 13602 8316
rect 13633 8313 13645 8316
rect 13679 8313 13691 8347
rect 13633 8307 13691 8313
rect 12158 8276 12164 8288
rect 11440 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 2222 8032 2228 8084
rect 2280 8032 2286 8084
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 3605 8075 3663 8081
rect 2731 8044 3096 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 2409 8007 2467 8013
rect 2409 7973 2421 8007
rect 2455 8004 2467 8007
rect 2455 7976 2774 8004
rect 2455 7973 2467 7976
rect 2409 7967 2467 7973
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 2406 7868 2412 7880
rect 2179 7840 2412 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2556 7840 2605 7868
rect 2556 7828 2562 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2746 7868 2774 7976
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2746 7840 2881 7868
rect 2593 7831 2651 7837
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 3068 7868 3096 8044
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 4154 8072 4160 8084
rect 3651 8044 4160 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4338 8032 4344 8084
rect 4396 8032 4402 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5040 8044 5181 8072
rect 5040 8032 5046 8044
rect 5169 8041 5181 8044
rect 5215 8072 5227 8075
rect 5215 8044 7043 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 4356 8004 4384 8032
rect 6914 8004 6920 8016
rect 3160 7976 4384 8004
rect 5368 7976 6920 8004
rect 3160 7945 3188 7976
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7905 3203 7939
rect 3878 7936 3884 7948
rect 3145 7899 3203 7905
rect 3252 7908 3884 7936
rect 3252 7868 3280 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4430 7896 4436 7948
rect 4488 7896 4494 7948
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4540 7908 4997 7936
rect 3068 7840 3280 7868
rect 2961 7831 3019 7837
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 2976 7800 3004 7831
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3476 7840 3801 7868
rect 3476 7828 3482 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4540 7868 4568 7908
rect 4985 7905 4997 7908
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 4120 7840 4568 7868
rect 4120 7828 4126 7840
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 5368 7877 5396 7976
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 7015 8004 7043 8044
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 8570 8072 8576 8084
rect 7156 8044 8576 8072
rect 7156 8032 7162 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 8904 8044 9229 8072
rect 8904 8032 8910 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 11882 8072 11888 8084
rect 9364 8044 11888 8072
rect 9364 8032 9370 8044
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 14148 8044 14197 8072
rect 14148 8032 14154 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 10042 8004 10048 8016
rect 7015 7976 10048 8004
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 6012 7908 6224 7936
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4672 7840 5089 7868
rect 4672 7828 4678 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5500 7840 5549 7868
rect 5500 7828 5506 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 6012 7809 6040 7908
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 2976 7772 6009 7800
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 1673 7735 1731 7741
rect 1673 7732 1685 7735
rect 1636 7704 1685 7732
rect 1636 7692 1642 7704
rect 1673 7701 1685 7704
rect 1719 7701 1731 7735
rect 1673 7695 1731 7701
rect 3878 7692 3884 7744
rect 3936 7692 3942 7744
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4706 7732 4712 7744
rect 4111 7704 4712 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 6104 7732 6132 7831
rect 6196 7800 6224 7908
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6696 7908 6837 7936
rect 6696 7896 6702 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 9214 7936 9220 7948
rect 7055 7908 9220 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 9950 7936 9956 7948
rect 9447 7908 9956 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13814 7936 13820 7948
rect 13127 7908 13820 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 7282 7868 7288 7880
rect 6319 7840 7288 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7650 7868 7656 7880
rect 7432 7840 7656 7868
rect 7432 7828 7438 7840
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8938 7868 8944 7880
rect 8343 7840 8944 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7868 9091 7871
rect 9122 7868 9128 7880
rect 9079 7840 9128 7868
rect 9079 7837 9091 7840
rect 9033 7831 9091 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 10045 7871 10103 7877
rect 10045 7868 10057 7871
rect 9640 7840 10057 7868
rect 9640 7828 9646 7840
rect 10045 7837 10057 7840
rect 10091 7868 10103 7871
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 10091 7840 11529 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 11517 7837 11529 7840
rect 11563 7868 11575 7871
rect 11606 7868 11612 7880
rect 11563 7840 11612 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 11784 7871 11842 7877
rect 11784 7837 11796 7871
rect 11830 7868 11842 7871
rect 12802 7868 12808 7880
rect 11830 7840 12808 7868
rect 11830 7837 11842 7840
rect 11784 7831 11842 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13964 7840 14105 7868
rect 13964 7828 13970 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 6733 7803 6791 7809
rect 6733 7800 6745 7803
rect 6196 7772 6745 7800
rect 6733 7769 6745 7772
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 7098 7760 7104 7812
rect 7156 7760 7162 7812
rect 7469 7803 7527 7809
rect 7469 7769 7481 7803
rect 7515 7800 7527 7803
rect 8478 7800 8484 7812
rect 7515 7772 8484 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 9953 7803 10011 7809
rect 8619 7772 9904 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 7116 7732 7144 7760
rect 6104 7704 7144 7732
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 7708 7704 8217 7732
rect 7708 7692 7714 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 8386 7692 8392 7744
rect 8444 7692 8450 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9398 7732 9404 7744
rect 8812 7704 9404 7732
rect 8812 7692 8818 7704
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 9876 7732 9904 7772
rect 9953 7769 9965 7803
rect 9999 7800 10011 7803
rect 10290 7803 10348 7809
rect 10290 7800 10302 7803
rect 9999 7772 10302 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 10290 7769 10302 7772
rect 10336 7769 10348 7803
rect 12710 7800 12716 7812
rect 10290 7763 10348 7769
rect 10520 7772 12716 7800
rect 10520 7732 10548 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7800 13231 7803
rect 13446 7800 13452 7812
rect 13219 7772 13452 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 13725 7803 13783 7809
rect 13725 7800 13737 7803
rect 13596 7772 13737 7800
rect 13596 7760 13602 7772
rect 13725 7769 13737 7772
rect 13771 7769 13783 7803
rect 13725 7763 13783 7769
rect 9876 7704 10548 7732
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11425 7735 11483 7741
rect 11425 7732 11437 7735
rect 11112 7704 11437 7732
rect 11112 7692 11118 7704
rect 11425 7701 11437 7704
rect 11471 7701 11483 7735
rect 11425 7695 11483 7701
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12802 7732 12808 7744
rect 12676 7704 12808 7732
rect 12676 7692 12682 7704
rect 12802 7692 12808 7704
rect 12860 7732 12866 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12860 7704 12909 7732
rect 12860 7692 12866 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 1949 7531 2007 7537
rect 1949 7497 1961 7531
rect 1995 7528 2007 7531
rect 2130 7528 2136 7540
rect 1995 7500 2136 7528
rect 1995 7497 2007 7500
rect 1949 7491 2007 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9582 7528 9588 7540
rect 9355 7500 9588 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10428 7500 13584 7528
rect 1872 7432 3096 7460
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 1872 7401 1900 7432
rect 3068 7404 3096 7432
rect 3326 7420 3332 7472
rect 3384 7420 3390 7472
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 3936 7432 4660 7460
rect 3936 7420 3942 7432
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 2332 7324 2360 7355
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 3050 7352 3056 7404
rect 3108 7352 3114 7404
rect 3344 7324 3372 7420
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4632 7401 4660 7432
rect 4706 7420 4712 7472
rect 4764 7420 4770 7472
rect 5718 7420 5724 7472
rect 5776 7460 5782 7472
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 5776 7432 6561 7460
rect 5776 7420 5782 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 6549 7423 6607 7429
rect 7282 7420 7288 7472
rect 7340 7420 7346 7472
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8202 7460 8208 7472
rect 7883 7432 8208 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 8404 7460 8432 7488
rect 10428 7460 10456 7500
rect 8404 7432 10456 7460
rect 11701 7463 11759 7469
rect 11701 7429 11713 7463
rect 11747 7460 11759 7463
rect 13446 7460 13452 7472
rect 11747 7432 13452 7460
rect 11747 7429 11759 7432
rect 11701 7423 11759 7429
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 4617 7395 4675 7401
rect 4028 7364 4568 7392
rect 4028 7352 4034 7364
rect 1452 7296 3372 7324
rect 4433 7327 4491 7333
rect 1452 7284 1458 7296
rect 4433 7293 4445 7327
rect 4479 7293 4491 7327
rect 4540 7324 4568 7364
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4724 7392 4752 7420
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4724 7364 5181 7392
rect 4617 7355 4675 7361
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5994 7352 6000 7404
rect 6052 7352 6058 7404
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7392 7392 7420 7420
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7392 7364 7665 7392
rect 7193 7355 7251 7361
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 9944 7395 10002 7401
rect 9944 7361 9956 7395
rect 9990 7392 10002 7395
rect 10226 7392 10232 7404
rect 9990 7364 10232 7392
rect 9990 7361 10002 7364
rect 9944 7355 10002 7361
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 4540 7296 5365 7324
rect 4433 7287 4491 7293
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 5353 7287 5411 7293
rect 5552 7296 6469 7324
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 3142 7256 3148 7268
rect 1627 7228 3148 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 3881 7259 3939 7265
rect 3881 7256 3893 7259
rect 3844 7228 3893 7256
rect 3844 7216 3850 7228
rect 3881 7225 3893 7228
rect 3927 7225 3939 7259
rect 3881 7219 3939 7225
rect 2406 7148 2412 7200
rect 2464 7148 2470 7200
rect 4448 7188 4476 7287
rect 4982 7216 4988 7268
rect 5040 7216 5046 7268
rect 5552 7265 5580 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 7208 7324 7236 7355
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 13556 7401 13584 7500
rect 13906 7488 13912 7540
rect 13964 7488 13970 7540
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 11072 7364 11345 7392
rect 6457 7287 6515 7293
rect 6564 7296 7236 7324
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5123 7228 5549 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5537 7225 5549 7228
rect 5583 7225 5595 7259
rect 5537 7219 5595 7225
rect 5994 7216 6000 7268
rect 6052 7256 6058 7268
rect 6564 7256 6592 7296
rect 8294 7284 8300 7336
rect 8352 7284 8358 7336
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 8444 7296 9689 7324
rect 8444 7284 8450 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 6052 7228 6592 7256
rect 7009 7259 7067 7265
rect 6052 7216 6058 7228
rect 7009 7225 7021 7259
rect 7055 7225 7067 7259
rect 7009 7219 7067 7225
rect 7469 7259 7527 7265
rect 7469 7225 7481 7259
rect 7515 7256 7527 7259
rect 8312 7256 8340 7284
rect 7515 7228 8340 7256
rect 7515 7225 7527 7228
rect 7469 7219 7527 7225
rect 5000 7188 5028 7216
rect 4448 7160 5028 7188
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 6012 7188 6040 7216
rect 5316 7160 6040 7188
rect 6089 7191 6147 7197
rect 5316 7148 5322 7160
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 6638 7188 6644 7200
rect 6135 7160 6644 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7024 7188 7052 7219
rect 7098 7188 7104 7200
rect 7024 7160 7104 7188
rect 7098 7148 7104 7160
rect 7156 7188 7162 7200
rect 8294 7188 8300 7200
rect 7156 7160 8300 7188
rect 7156 7148 7162 7160
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10962 7188 10968 7200
rect 10008 7160 10968 7188
rect 10008 7148 10014 7160
rect 10962 7148 10968 7160
rect 11020 7188 11026 7200
rect 11072 7197 11100 7364
rect 11333 7361 11345 7364
rect 11379 7361 11391 7395
rect 11333 7355 11391 7361
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13924 7392 13952 7488
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13924 7364 14289 7392
rect 13541 7355 13599 7361
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7324 11667 7327
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 11655 7296 12357 7324
rect 11655 7293 11667 7296
rect 11609 7287 11667 7293
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 12802 7324 12808 7336
rect 12759 7296 12808 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 11698 7216 11704 7268
rect 11756 7256 11762 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 11756 7228 12173 7256
rect 11756 7216 11762 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 13372 7256 13400 7287
rect 12161 7219 12219 7225
rect 12406 7228 13400 7256
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 11020 7160 11069 7188
rect 11020 7148 11026 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 12406 7188 12434 7228
rect 11940 7160 12434 7188
rect 11940 7148 11946 7160
rect 13262 7148 13268 7200
rect 13320 7148 13326 7200
rect 13906 7148 13912 7200
rect 13964 7148 13970 7200
rect 14090 7148 14096 7200
rect 14148 7148 14154 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3513 6987 3571 6993
rect 3513 6984 3525 6987
rect 3108 6956 3525 6984
rect 3108 6944 3114 6956
rect 3513 6953 3525 6956
rect 3559 6984 3571 6987
rect 5258 6984 5264 6996
rect 3559 6956 5264 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5442 6944 5448 6996
rect 5500 6944 5506 6996
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 6178 6984 6184 6996
rect 5684 6956 6184 6984
rect 5684 6944 5690 6956
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 7006 6984 7012 6996
rect 6604 6956 7012 6984
rect 6604 6944 6610 6956
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 8938 6944 8944 6996
rect 8996 6944 9002 6996
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 11606 6984 11612 6996
rect 9548 6956 11612 6984
rect 9548 6944 9554 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 13449 6987 13507 6993
rect 13449 6953 13461 6987
rect 13495 6984 13507 6987
rect 14274 6984 14280 6996
rect 13495 6956 14280 6984
rect 13495 6953 13507 6956
rect 13449 6947 13507 6953
rect 6365 6919 6423 6925
rect 4908 6888 5941 6916
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 2774 6780 2780 6792
rect 2179 6752 2780 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 2832 6752 3801 6780
rect 2832 6740 2838 6752
rect 3789 6749 3801 6752
rect 3835 6780 3847 6783
rect 3878 6780 3884 6792
rect 3835 6752 3884 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4062 6789 4068 6792
rect 4056 6780 4068 6789
rect 4023 6752 4068 6780
rect 4056 6743 4068 6752
rect 4062 6740 4068 6743
rect 4120 6740 4126 6792
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6712 2099 6715
rect 2378 6715 2436 6721
rect 2378 6712 2390 6715
rect 2087 6684 2390 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 2378 6681 2390 6684
rect 2424 6681 2436 6715
rect 2378 6675 2436 6681
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 4908 6644 4936 6888
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5040 6820 5825 6848
rect 5040 6808 5046 6820
rect 5813 6817 5825 6820
rect 5859 6817 5871 6851
rect 5913 6848 5941 6888
rect 6365 6885 6377 6919
rect 6411 6916 6423 6919
rect 7098 6916 7104 6928
rect 6411 6888 7104 6916
rect 6411 6885 6423 6888
rect 6365 6879 6423 6885
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 8956 6916 8984 6944
rect 8956 6888 12112 6916
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 5913 6820 6561 6848
rect 5813 6811 5871 6817
rect 6549 6817 6561 6820
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 8864 6820 9904 6848
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5629 6783 5687 6789
rect 5629 6780 5641 6783
rect 5500 6752 5641 6780
rect 5500 6740 5506 6752
rect 5629 6749 5641 6752
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 8386 6780 8392 6792
rect 7423 6752 8392 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 7650 6721 7656 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5736 6684 5917 6712
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 3476 6616 5181 6644
rect 3476 6604 3482 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5736 6644 5764 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 7644 6712 7656 6721
rect 7611 6684 7656 6712
rect 5905 6675 5963 6681
rect 7644 6675 7656 6684
rect 7650 6672 7656 6675
rect 7708 6672 7714 6724
rect 5316 6616 5764 6644
rect 5316 6604 5322 6616
rect 7190 6604 7196 6656
rect 7248 6604 7254 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 8864 6644 8892 6820
rect 9876 6789 9904 6820
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 11241 6851 11299 6857
rect 10468 6820 10640 6848
rect 10468 6808 10474 6820
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 9907 6752 10517 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 9033 6715 9091 6721
rect 9033 6712 9045 6715
rect 8956 6684 9045 6712
rect 8956 6656 8984 6684
rect 9033 6681 9045 6684
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 9125 6715 9183 6721
rect 9125 6681 9137 6715
rect 9171 6681 9183 6715
rect 9125 6675 9183 6681
rect 8812 6616 8892 6644
rect 8812 6604 8818 6616
rect 8938 6604 8944 6656
rect 8996 6604 9002 6656
rect 9140 6644 9168 6675
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 9677 6715 9735 6721
rect 9677 6712 9689 6715
rect 9272 6684 9689 6712
rect 9272 6672 9278 6684
rect 9677 6681 9689 6684
rect 9723 6681 9735 6715
rect 9677 6675 9735 6681
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 10413 6715 10471 6721
rect 10413 6712 10425 6715
rect 10284 6684 10425 6712
rect 10284 6672 10290 6684
rect 10413 6681 10425 6684
rect 10459 6681 10471 6715
rect 10612 6712 10640 6820
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11606 6848 11612 6860
rect 11287 6820 11612 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 11882 6808 11888 6860
rect 11940 6808 11946 6860
rect 12084 6848 12112 6888
rect 12084 6820 12204 6848
rect 11900 6780 11928 6808
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11900 6752 12081 6780
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 10612 6684 11345 6712
rect 10413 6675 10471 6681
rect 11333 6681 11345 6684
rect 11379 6681 11391 6715
rect 11333 6675 11391 6681
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 11885 6715 11943 6721
rect 11885 6712 11897 6715
rect 11756 6684 11897 6712
rect 11756 6672 11762 6684
rect 11885 6681 11897 6684
rect 11931 6681 11943 6715
rect 12176 6712 12204 6820
rect 12336 6783 12394 6789
rect 12336 6749 12348 6783
rect 12382 6780 12394 6783
rect 13262 6780 13268 6792
rect 12382 6752 13268 6780
rect 12382 6749 12394 6752
rect 12336 6743 12394 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 12176 6684 12434 6712
rect 11885 6675 11943 6681
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 9140 6616 10609 6644
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10597 6607 10655 6613
rect 10778 6604 10784 6656
rect 10836 6604 10842 6656
rect 12406 6644 12434 6684
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 13078 6712 13084 6724
rect 12676 6684 13084 6712
rect 12676 6672 12682 6684
rect 13078 6672 13084 6684
rect 13136 6672 13142 6724
rect 13464 6644 13492 6947
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 13722 6916 13728 6928
rect 13596 6888 13728 6916
rect 13596 6876 13602 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13872 6820 14105 6848
rect 13872 6808 13878 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 13538 6740 13544 6792
rect 13596 6740 13602 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13998 6780 14004 6792
rect 13679 6752 14004 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 13814 6644 13820 6656
rect 12406 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 3881 6443 3939 6449
rect 2464 6412 3188 6440
rect 2464 6400 2470 6412
rect 3160 6381 3188 6412
rect 3881 6409 3893 6443
rect 3927 6440 3939 6443
rect 3970 6440 3976 6452
rect 3927 6412 3976 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 5132 6412 5549 6440
rect 5132 6400 5138 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5810 6440 5816 6452
rect 5537 6403 5595 6409
rect 5736 6412 5816 6440
rect 3145 6375 3203 6381
rect 1412 6344 2774 6372
rect 1412 6313 1440 6344
rect 2746 6316 2774 6344
rect 3145 6341 3157 6375
rect 3191 6341 3203 6375
rect 3145 6335 3203 6341
rect 4424 6375 4482 6381
rect 4424 6341 4436 6375
rect 4470 6372 4482 6375
rect 5552 6372 5580 6403
rect 5736 6372 5764 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5960 6412 6193 6440
rect 5960 6400 5966 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 7742 6440 7748 6452
rect 7432 6412 7748 6440
rect 7432 6400 7438 6412
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8478 6440 8484 6452
rect 8343 6412 8484 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9079 6412 9536 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 7190 6372 7196 6384
rect 4470 6344 5404 6372
rect 5552 6344 5764 6372
rect 5828 6344 7196 6372
rect 4470 6341 4482 6344
rect 4424 6335 4482 6341
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1664 6307 1722 6313
rect 1664 6273 1676 6307
rect 1710 6304 1722 6307
rect 2222 6304 2228 6316
rect 1710 6276 2228 6304
rect 1710 6273 1722 6276
rect 1664 6267 1722 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2746 6276 2780 6316
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3752 6276 4077 6304
rect 3752 6264 3758 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 5376 6304 5404 6344
rect 5828 6304 5856 6344
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 4856 6276 5212 6304
rect 5376 6276 5856 6304
rect 4856 6264 4862 6276
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3099 6208 3832 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3326 6128 3332 6180
rect 3384 6128 3390 6180
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6137 3663 6171
rect 3804 6168 3832 6208
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 3936 6208 4169 6236
rect 3936 6196 3942 6208
rect 3970 6168 3976 6180
rect 3804 6140 3976 6168
rect 3605 6131 3663 6137
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 3344 6100 3372 6128
rect 2823 6072 3372 6100
rect 3620 6100 3648 6131
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4080 6112 4108 6208
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 5184 6168 5212 6276
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6043 6276 7113 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5500 6208 5764 6236
rect 5500 6196 5506 6208
rect 5626 6168 5632 6180
rect 5184 6140 5632 6168
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 5736 6177 5764 6208
rect 5721 6171 5779 6177
rect 5721 6137 5733 6171
rect 5767 6137 5779 6171
rect 5721 6131 5779 6137
rect 3878 6100 3884 6112
rect 3620 6072 3884 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4062 6060 4068 6112
rect 4120 6060 4126 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 6012 6100 6040 6267
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7432 6276 7573 6304
rect 7432 6264 7438 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6144 6208 6469 6236
rect 6144 6196 6150 6208
rect 6457 6205 6469 6208
rect 6503 6236 6515 6239
rect 6914 6236 6920 6248
rect 6503 6208 6920 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 7064 6208 7205 6236
rect 7064 6196 7070 6208
rect 7193 6205 7205 6208
rect 7239 6236 7251 6239
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 7239 6208 7665 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7653 6205 7665 6208
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 7834 6196 7840 6248
rect 7892 6196 7898 6248
rect 8496 6236 8524 6400
rect 8588 6372 8616 6403
rect 9508 6381 9536 6412
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 10962 6400 10968 6452
rect 11020 6400 11026 6452
rect 11698 6440 11704 6452
rect 11256 6412 11704 6440
rect 9493 6375 9551 6381
rect 8588 6344 9260 6372
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 9232 6313 9260 6344
rect 9493 6341 9505 6375
rect 9539 6341 9551 6375
rect 9876 6372 9904 6400
rect 10873 6375 10931 6381
rect 10873 6372 10885 6375
rect 9876 6344 10885 6372
rect 9493 6335 9551 6341
rect 10873 6341 10885 6344
rect 10919 6341 10931 6375
rect 10873 6335 10931 6341
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 10778 6304 10784 6316
rect 9217 6267 9275 6273
rect 10060 6276 10784 6304
rect 8938 6236 8944 6248
rect 8496 6208 8944 6236
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 6178 6128 6184 6180
rect 6236 6168 6242 6180
rect 9140 6168 9168 6264
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6236 9459 6239
rect 10060 6236 10088 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10980 6313 11008 6400
rect 11256 6384 11284 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 13538 6440 13544 6452
rect 11799 6412 13544 6440
rect 11238 6332 11244 6384
rect 11296 6332 11302 6384
rect 11799 6372 11827 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 14366 6400 14372 6452
rect 14424 6400 14430 6452
rect 11624 6344 11827 6372
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 9447 6208 10088 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 10134 6196 10140 6248
rect 10192 6236 10198 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10192 6208 10241 6236
rect 10192 6196 10198 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 11624 6236 11652 6344
rect 12802 6332 12808 6384
rect 12860 6372 12866 6384
rect 12860 6344 14320 6372
rect 12860 6332 12866 6344
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 14292 6313 14320 6344
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 12336 6307 12394 6313
rect 12336 6273 12348 6307
rect 12382 6304 12394 6307
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 12382 6276 14197 6304
rect 12382 6273 12394 6276
rect 12336 6267 12394 6273
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 11808 6236 11836 6267
rect 10229 6199 10287 6205
rect 10888 6208 11652 6236
rect 11716 6208 11836 6236
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 6236 6140 7420 6168
rect 9140 6140 9965 6168
rect 6236 6128 6242 6140
rect 4396 6072 6040 6100
rect 4396 6060 4402 6072
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 7392 6109 7420 6140
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 10686 6168 10692 6180
rect 10560 6140 10692 6168
rect 10560 6128 10566 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6144 6072 7021 6100
rect 6144 6060 6150 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6069 7435 6103
rect 7377 6063 7435 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 10888 6100 10916 6208
rect 11716 6180 11744 6208
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11940 6208 12081 6236
rect 11940 6196 11946 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 13814 6236 13820 6248
rect 13679 6208 13820 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11020 6140 11529 6168
rect 11020 6128 11026 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 11698 6128 11704 6180
rect 11756 6128 11762 6180
rect 13096 6168 13124 6196
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 13096 6140 13461 6168
rect 13449 6137 13461 6140
rect 13495 6137 13507 6171
rect 13449 6131 13507 6137
rect 8352 6072 10916 6100
rect 8352 6060 8358 6072
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11480 6072 11897 6100
rect 11480 6060 11486 6072
rect 11885 6069 11897 6072
rect 11931 6069 11943 6103
rect 11885 6063 11943 6069
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 13998 6100 14004 6112
rect 12308 6072 14004 6100
rect 12308 6060 12314 6072
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1762 5896 1768 5908
rect 1627 5868 1768 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 3050 5856 3056 5908
rect 3108 5856 3114 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3694 5896 3700 5908
rect 3467 5868 3700 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3844 5868 3985 5896
rect 3844 5856 3850 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 5258 5896 5264 5908
rect 4663 5868 5264 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6457 5899 6515 5905
rect 6457 5896 6469 5899
rect 6052 5868 6469 5896
rect 6052 5856 6058 5868
rect 6457 5865 6469 5868
rect 6503 5896 6515 5899
rect 6730 5896 6736 5908
rect 6503 5868 6736 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7190 5856 7196 5908
rect 7248 5856 7254 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 7524 5868 7573 5896
rect 7524 5856 7530 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7892 5868 8033 5896
rect 7892 5856 7898 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8435 5868 10548 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 3068 5828 3096 5856
rect 1780 5800 3096 5828
rect 3237 5831 3295 5837
rect 1780 5701 1808 5800
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 3878 5828 3884 5840
rect 3283 5800 3884 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 3878 5788 3884 5800
rect 3936 5828 3942 5840
rect 4706 5828 4712 5840
rect 3936 5800 4712 5828
rect 3936 5788 3942 5800
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 4798 5788 4804 5840
rect 4856 5788 4862 5840
rect 5074 5828 5080 5840
rect 4908 5800 5080 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 1946 5760 1952 5772
rect 1903 5732 1952 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 2038 5720 2044 5772
rect 2096 5720 2102 5772
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3418 5760 3424 5772
rect 2740 5732 3424 5760
rect 2740 5720 2746 5732
rect 3418 5720 3424 5732
rect 3476 5760 3482 5772
rect 3476 5732 3648 5760
rect 3476 5720 3482 5732
rect 3620 5701 3648 5732
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3651 5664 4169 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4908 5692 4936 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 6638 5788 6644 5840
rect 6696 5788 6702 5840
rect 7374 5828 7380 5840
rect 7116 5800 7380 5828
rect 5000 5732 5212 5760
rect 5000 5701 5028 5732
rect 4571 5664 4936 5692
rect 4985 5695 5043 5701
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 1946 5584 1952 5636
rect 2004 5624 2010 5636
rect 2222 5624 2228 5636
rect 2004 5596 2228 5624
rect 2004 5584 2010 5596
rect 2222 5584 2228 5596
rect 2280 5584 2286 5636
rect 2406 5584 2412 5636
rect 2464 5624 2470 5636
rect 2501 5627 2559 5633
rect 2501 5624 2513 5627
rect 2464 5596 2513 5624
rect 2464 5584 2470 5596
rect 2501 5593 2513 5596
rect 2547 5624 2559 5627
rect 2685 5627 2743 5633
rect 2685 5624 2697 5627
rect 2547 5596 2697 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 2685 5593 2697 5596
rect 2731 5593 2743 5627
rect 2685 5587 2743 5593
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5593 2835 5627
rect 5092 5624 5120 5655
rect 2777 5587 2835 5593
rect 5000 5596 5120 5624
rect 5184 5624 5212 5732
rect 5344 5695 5402 5701
rect 5344 5661 5356 5695
rect 5390 5692 5402 5695
rect 5902 5692 5908 5704
rect 5390 5664 5908 5692
rect 5390 5661 5402 5664
rect 5344 5655 5402 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6656 5701 6684 5788
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7116 5692 7144 5800
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 8754 5828 8760 5840
rect 8312 5800 8760 5828
rect 7208 5732 7696 5760
rect 7208 5704 7236 5732
rect 7064 5664 7144 5692
rect 7064 5652 7070 5664
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7668 5701 7696 5732
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 5626 5624 5632 5636
rect 5184 5596 5632 5624
rect 2792 5556 2820 5587
rect 5000 5568 5028 5596
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 7392 5624 7420 5655
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8312 5701 8340 5800
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10321 5831 10379 5837
rect 10321 5828 10333 5831
rect 10192 5800 10333 5828
rect 10192 5788 10198 5800
rect 10321 5797 10333 5800
rect 10367 5797 10379 5831
rect 10321 5791 10379 5797
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8404 5732 8953 5760
rect 8404 5704 8432 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10100 5732 10425 5760
rect 10100 5720 10106 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7800 5664 7941 5692
rect 7800 5652 7806 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 8588 5624 8616 5655
rect 6144 5596 7420 5624
rect 7484 5596 8616 5624
rect 9208 5627 9266 5633
rect 6144 5584 6150 5596
rect 3418 5556 3424 5568
rect 2792 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 4341 5559 4399 5565
rect 4341 5556 4353 5559
rect 3936 5528 4353 5556
rect 3936 5516 3942 5528
rect 4341 5525 4353 5528
rect 4387 5525 4399 5559
rect 4341 5519 4399 5525
rect 4982 5516 4988 5568
rect 5040 5516 5046 5568
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 7484 5556 7512 5596
rect 9208 5593 9220 5627
rect 9254 5624 9266 5627
rect 9858 5624 9864 5636
rect 9254 5596 9864 5624
rect 9254 5593 9266 5596
rect 9208 5587 9266 5593
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 5316 5528 7512 5556
rect 5316 5516 5322 5528
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7708 5528 7757 5556
rect 7708 5516 7714 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 8665 5559 8723 5565
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 10410 5556 10416 5568
rect 8711 5528 10416 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10520 5556 10548 5868
rect 10962 5856 10968 5908
rect 11020 5856 11026 5908
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 11422 5856 11428 5908
rect 11480 5856 11486 5908
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 12250 5856 12256 5908
rect 12308 5856 12314 5908
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13504 5868 14105 5896
rect 13504 5856 13510 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10980 5760 11008 5856
rect 10643 5732 11008 5760
rect 11072 5760 11100 5856
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11072 5732 11345 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 11020 5664 11161 5692
rect 11020 5652 11026 5664
rect 11149 5661 11161 5664
rect 11195 5692 11207 5695
rect 11440 5692 11468 5856
rect 11195 5664 11468 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 11057 5627 11115 5633
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 11624 5624 11652 5856
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 11974 5760 11980 5772
rect 11931 5732 11980 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 11103 5596 11652 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 12084 5624 12112 5655
rect 12032 5596 12112 5624
rect 12032 5584 12038 5596
rect 12268 5556 12296 5856
rect 13906 5828 13912 5840
rect 13280 5800 13912 5828
rect 13280 5769 13308 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12676 5664 12725 5692
rect 12676 5652 12682 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 12342 5584 12348 5636
rect 12400 5624 12406 5636
rect 13357 5627 13415 5633
rect 12400 5596 12664 5624
rect 12400 5584 12406 5596
rect 10520 5528 12296 5556
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 12492 5528 12541 5556
rect 12492 5516 12498 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12636 5556 12664 5596
rect 13357 5593 13369 5627
rect 13403 5593 13415 5627
rect 13357 5587 13415 5593
rect 13909 5627 13967 5633
rect 13909 5593 13921 5627
rect 13955 5624 13967 5627
rect 14366 5624 14372 5636
rect 13955 5596 14372 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12636 5528 12817 5556
rect 12529 5519 12587 5525
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 13372 5556 13400 5587
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 14550 5556 14556 5568
rect 13372 5528 14556 5556
rect 12805 5519 12863 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1360 5324 1440 5352
rect 1360 5312 1366 5324
rect 1412 5216 1440 5324
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 2004 5324 2237 5352
rect 2004 5312 2010 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 4246 5352 4252 5364
rect 3108 5324 4252 5352
rect 3108 5312 3114 5324
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5132 5324 5825 5352
rect 5132 5312 5138 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 6362 5352 6368 5364
rect 5813 5315 5871 5321
rect 5920 5324 6368 5352
rect 1762 5244 1768 5296
rect 1820 5284 1826 5296
rect 2409 5287 2467 5293
rect 2409 5284 2421 5287
rect 1820 5256 2421 5284
rect 1820 5244 1826 5256
rect 2409 5253 2421 5256
rect 2455 5253 2467 5287
rect 2409 5247 2467 5253
rect 2498 5244 2504 5296
rect 2556 5284 2562 5296
rect 2593 5287 2651 5293
rect 2593 5284 2605 5287
rect 2556 5256 2605 5284
rect 2556 5244 2562 5256
rect 2593 5253 2605 5256
rect 2639 5284 2651 5287
rect 2639 5256 5856 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 5828 5228 5856 5256
rect 2222 5216 2228 5228
rect 1412 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 4120 5188 4353 5216
rect 4120 5176 4126 5188
rect 4341 5185 4353 5188
rect 4387 5216 4399 5219
rect 4982 5216 4988 5228
rect 4387 5188 4988 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5534 5216 5540 5228
rect 5215 5188 5540 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5810 5176 5816 5228
rect 5868 5176 5874 5228
rect 5920 5216 5948 5324
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 6696 5324 6745 5352
rect 6696 5312 6702 5324
rect 6733 5321 6745 5324
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 6880 5324 7389 5352
rect 6880 5312 6886 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 9950 5352 9956 5364
rect 7377 5315 7435 5321
rect 7760 5324 9956 5352
rect 6089 5287 6147 5293
rect 6089 5253 6101 5287
rect 6135 5284 6147 5287
rect 7760 5284 7788 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10962 5352 10968 5364
rect 10428 5324 10968 5352
rect 6135 5256 7788 5284
rect 7837 5287 7895 5293
rect 6135 5253 6147 5256
rect 6089 5247 6147 5253
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8202 5284 8208 5296
rect 7883 5256 8208 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 10428 5293 10456 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12066 5352 12072 5364
rect 11931 5324 12072 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 14090 5312 14096 5364
rect 14148 5312 14154 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14240 5324 14289 5352
rect 14240 5312 14246 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 10413 5287 10471 5293
rect 8312 5256 9812 5284
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5920 5188 6009 5216
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6236 5188 6561 5216
rect 6236 5176 6242 5188
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 6822 5216 6828 5228
rect 6595 5188 6828 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6972 5188 7021 5216
rect 6972 5176 6978 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 3326 5148 3332 5160
rect 1719 5120 3332 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 3326 5108 3332 5120
rect 3384 5148 3390 5160
rect 3602 5148 3608 5160
rect 3384 5120 3608 5148
rect 3384 5108 3390 5120
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 4212 5120 4445 5148
rect 4212 5108 4218 5120
rect 4433 5117 4445 5120
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 1762 5040 1768 5092
rect 1820 5080 1826 5092
rect 4632 5080 4660 5111
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5626 5108 5632 5160
rect 5684 5108 5690 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 7576 5148 7604 5179
rect 5960 5120 7604 5148
rect 5960 5108 5966 5120
rect 1820 5052 4660 5080
rect 5644 5080 5672 5108
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 5644 5052 6837 5080
rect 1820 5040 1826 5052
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 8312 5080 8340 5256
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 6825 5043 6883 5049
rect 7116 5052 8340 5080
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 7116 5012 7144 5052
rect 8386 5040 8392 5092
rect 8444 5080 8450 5092
rect 9214 5080 9220 5092
rect 8444 5052 9220 5080
rect 8444 5040 8450 5052
rect 9214 5040 9220 5052
rect 9272 5080 9278 5092
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 9272 5052 9321 5080
rect 9272 5040 9278 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9692 5080 9720 5179
rect 9784 5148 9812 5256
rect 10413 5253 10425 5287
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 10505 5287 10563 5293
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 12618 5284 12624 5296
rect 10551 5256 12624 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 12710 5244 12716 5296
rect 12768 5284 12774 5296
rect 13541 5287 13599 5293
rect 13541 5284 13553 5287
rect 12768 5256 13553 5284
rect 12768 5244 12774 5256
rect 13541 5253 13553 5256
rect 13587 5253 13599 5287
rect 13541 5247 13599 5253
rect 13630 5244 13636 5296
rect 13688 5244 13694 5296
rect 14108 5284 14136 5312
rect 14108 5256 14504 5284
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10042 5216 10048 5228
rect 9999 5188 10048 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11606 5216 11612 5228
rect 11379 5188 11612 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 12244 5219 12302 5225
rect 12244 5185 12256 5219
rect 12290 5216 12302 5219
rect 13354 5216 13360 5228
rect 12290 5188 13360 5216
rect 12290 5185 12302 5188
rect 12244 5179 12302 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14476 5225 14504 5256
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 9784 5120 10701 5148
rect 10689 5117 10701 5120
rect 10735 5148 10747 5151
rect 11238 5148 11244 5160
rect 10735 5120 11244 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 11054 5080 11060 5092
rect 9692 5052 11060 5080
rect 9309 5043 9367 5049
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11716 5080 11744 5176
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11940 5120 11989 5148
rect 11940 5108 11946 5120
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 14093 5083 14151 5089
rect 11716 5052 11928 5080
rect 3844 4984 7144 5012
rect 7193 5015 7251 5021
rect 3844 4972 3850 4984
rect 7193 4981 7205 5015
rect 7239 5012 7251 5015
rect 8294 5012 8300 5024
rect 7239 4984 8300 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 9950 5012 9956 5024
rect 9815 4984 9956 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10042 4972 10048 5024
rect 10100 4972 10106 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11790 5012 11796 5024
rect 11195 4984 11796 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 11900 5012 11928 5052
rect 12912 5052 14044 5080
rect 12912 5012 12940 5052
rect 11900 4984 12940 5012
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13446 5012 13452 5024
rect 13403 4984 13452 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14016 5012 14044 5052
rect 14093 5049 14105 5083
rect 14139 5080 14151 5083
rect 14366 5080 14372 5092
rect 14139 5052 14372 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 14182 5012 14188 5024
rect 14016 4984 14188 5012
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 1228 4780 2360 4808
rect 1228 4752 1256 4780
rect 1210 4700 1216 4752
rect 1268 4700 1274 4752
rect 2332 4740 2360 4780
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2464 4780 3249 4808
rect 2464 4768 2470 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3878 4808 3884 4820
rect 3568 4780 3884 4808
rect 3568 4768 3574 4780
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4798 4808 4804 4820
rect 4304 4780 4804 4808
rect 4304 4768 4310 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6086 4808 6092 4820
rect 5960 4780 6092 4808
rect 5960 4768 5966 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 6880 4780 9674 4808
rect 6880 4768 6886 4780
rect 2332 4712 3096 4740
rect 3068 4681 3096 4712
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 3973 4743 4031 4749
rect 3973 4740 3985 4743
rect 3200 4712 3985 4740
rect 3200 4700 3206 4712
rect 3973 4709 3985 4712
rect 4019 4709 4031 4743
rect 3973 4703 4031 4709
rect 4157 4743 4215 4749
rect 4157 4709 4169 4743
rect 4203 4709 4215 4743
rect 4157 4703 4215 4709
rect 3053 4675 3111 4681
rect 2746 4644 3004 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 2746 4604 2774 4644
rect 1443 4576 2774 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 2866 4564 2872 4616
rect 2924 4564 2930 4616
rect 2976 4604 3004 4644
rect 3053 4641 3065 4675
rect 3099 4641 3111 4675
rect 4172 4672 4200 4703
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 5132 4712 6960 4740
rect 5132 4700 5138 4712
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 3053 4635 3111 4641
rect 3712 4644 4108 4672
rect 4172 4644 6837 4672
rect 3712 4604 3740 4644
rect 4080 4616 4108 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 6825 4635 6883 4641
rect 2976 4576 3740 4604
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 3970 4604 3976 4616
rect 3835 4576 3976 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 4304 4576 4353 4604
rect 4304 4564 4310 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4604 4675 4607
rect 4890 4604 4896 4616
rect 4663 4576 4896 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 1664 4539 1722 4545
rect 1664 4505 1676 4539
rect 1710 4536 1722 4539
rect 1710 4508 3648 4536
rect 1710 4505 1722 4508
rect 1664 4499 1722 4505
rect 2777 4471 2835 4477
rect 2777 4437 2789 4471
rect 2823 4468 2835 4471
rect 3326 4468 3332 4480
rect 2823 4440 3332 4468
rect 2823 4437 2835 4440
rect 2777 4431 2835 4437
rect 3326 4428 3332 4440
rect 3384 4428 3390 4480
rect 3620 4468 3648 4508
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 4448 4536 4476 4567
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 5132 4576 5181 4604
rect 5132 4564 5138 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 6932 4604 6960 4712
rect 9030 4700 9036 4752
rect 9088 4740 9094 4752
rect 9309 4743 9367 4749
rect 9309 4740 9321 4743
rect 9088 4712 9321 4740
rect 9088 4700 9094 4712
rect 9309 4709 9321 4712
rect 9355 4709 9367 4743
rect 9646 4740 9674 4780
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 9916 4780 10333 4808
rect 9916 4768 9922 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 10321 4771 10379 4777
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10652 4780 10885 4808
rect 10652 4768 10658 4780
rect 10873 4777 10885 4780
rect 10919 4808 10931 4811
rect 10962 4808 10968 4820
rect 10919 4780 10968 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11238 4768 11244 4820
rect 11296 4768 11302 4820
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 12434 4808 12440 4820
rect 11839 4780 12440 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13354 4768 13360 4820
rect 13412 4768 13418 4820
rect 13722 4808 13728 4820
rect 13464 4780 13728 4808
rect 10505 4743 10563 4749
rect 10505 4740 10517 4743
rect 9646 4712 10517 4740
rect 9309 4703 9367 4709
rect 10505 4709 10517 4712
rect 10551 4709 10563 4743
rect 11256 4740 11284 4768
rect 12529 4743 12587 4749
rect 12529 4740 12541 4743
rect 11256 4712 12541 4740
rect 10505 4703 10563 4709
rect 12529 4709 12541 4712
rect 12575 4709 12587 4743
rect 12529 4703 12587 4709
rect 8386 4632 8392 4684
rect 8444 4632 8450 4684
rect 8570 4632 8576 4684
rect 8628 4672 8634 4684
rect 9858 4672 9864 4684
rect 8628 4644 9864 4672
rect 8628 4632 8634 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10284 4644 10548 4672
rect 10284 4632 10290 4644
rect 6687 4576 6960 4604
rect 7377 4607 7435 4613
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 8404 4604 8432 4632
rect 7423 4576 8432 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 8938 4564 8944 4616
rect 8996 4564 9002 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 7006 4536 7012 4548
rect 3752 4508 4476 4536
rect 5000 4508 7012 4536
rect 3752 4496 3758 4508
rect 5000 4468 5028 4508
rect 7006 4496 7012 4508
rect 7064 4496 7070 4548
rect 7644 4539 7702 4545
rect 7644 4505 7656 4539
rect 7690 4536 7702 4539
rect 8386 4536 8392 4548
rect 7690 4508 8392 4536
rect 7690 4505 7702 4508
rect 7644 4499 7702 4505
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 9140 4536 9168 4567
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9272 4576 9689 4604
rect 9272 4564 9278 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 8496 4508 9168 4536
rect 3620 4440 5028 4468
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 5868 4440 6561 4468
rect 5868 4428 5874 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 7282 4428 7288 4480
rect 7340 4428 7346 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8496 4468 8524 4508
rect 7524 4440 8524 4468
rect 8757 4471 8815 4477
rect 7524 4428 7530 4440
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9232 4468 9260 4564
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10428 4536 10456 4567
rect 9548 4508 10456 4536
rect 9548 4496 9554 4508
rect 8803 4440 9260 4468
rect 10520 4468 10548 4644
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 11977 4675 12035 4681
rect 10652 4644 11376 4672
rect 10652 4632 10658 4644
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11348 4613 11376 4644
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12066 4672 12072 4684
rect 12023 4644 12072 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12802 4632 12808 4684
rect 12860 4632 12866 4684
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 11020 4576 11161 4604
rect 11020 4564 11026 4576
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11974 4496 11980 4548
rect 12032 4536 12038 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 12032 4508 12081 4536
rect 12032 4496 12038 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 13464 4536 13492 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13688 4576 14289 4604
rect 13688 4564 13694 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 12069 4499 12127 4505
rect 12406 4508 13492 4536
rect 12406 4468 12434 4508
rect 13538 4496 13544 4548
rect 13596 4496 13602 4548
rect 14369 4539 14427 4545
rect 14369 4536 14381 4539
rect 13648 4508 14381 4536
rect 10520 4440 12434 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 13648 4468 13676 4508
rect 14369 4505 14381 4508
rect 14415 4505 14427 4539
rect 14369 4499 14427 4505
rect 13504 4440 13676 4468
rect 13504 4428 13510 4440
rect 13814 4428 13820 4480
rect 13872 4428 13878 4480
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 1762 4224 1768 4276
rect 1820 4224 1826 4276
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 2280 4236 3648 4264
rect 2280 4224 2286 4236
rect 2498 4196 2504 4208
rect 1688 4168 2504 4196
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1578 4128 1584 4140
rect 1443 4100 1584 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 1688 4137 1716 4168
rect 2498 4156 2504 4168
rect 2556 4156 2562 4208
rect 3620 4196 3648 4236
rect 3694 4224 3700 4276
rect 3752 4224 3758 4276
rect 4433 4267 4491 4273
rect 4433 4233 4445 4267
rect 4479 4264 4491 4267
rect 4798 4264 4804 4276
rect 4479 4236 4804 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 5592 4236 5641 4264
rect 5592 4224 5598 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 6086 4264 6092 4276
rect 5767 4236 6092 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6420 4236 6960 4264
rect 6420 4224 6426 4236
rect 4338 4196 4344 4208
rect 3620 4168 4344 4196
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 6822 4196 6828 4208
rect 5828 4168 6828 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2958 4128 2964 4140
rect 2271 4100 2964 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 1026 4020 1032 4072
rect 1084 4060 1090 4072
rect 2148 4060 2176 4091
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3510 4128 3516 4140
rect 3099 4100 3516 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4632 4100 4905 4128
rect 1084 4032 2176 4060
rect 1084 4020 1090 4032
rect 2406 4020 2412 4072
rect 2464 4020 2470 4072
rect 2792 4032 3188 4060
rect 1489 3995 1547 4001
rect 1489 3961 1501 3995
rect 1535 3992 1547 3995
rect 2792 3992 2820 4032
rect 1535 3964 2820 3992
rect 3160 3992 3188 4032
rect 3234 4020 3240 4072
rect 3292 4020 3298 4072
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3384 4032 3985 4060
rect 3384 4020 3390 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 4632 4004 4660 4100
rect 4893 4097 4905 4100
rect 4939 4128 4951 4131
rect 5169 4131 5227 4137
rect 4939 4100 5120 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4856 4032 4997 4060
rect 4856 4020 4862 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 5092 4060 5120 4100
rect 5169 4097 5181 4131
rect 5215 4126 5227 4131
rect 5828 4128 5856 4168
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 6932 4196 6960 4236
rect 7006 4224 7012 4276
rect 7064 4224 7070 4276
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 8294 4224 8300 4276
rect 8352 4224 8358 4276
rect 8386 4224 8392 4276
rect 8444 4224 8450 4276
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 9030 4264 9036 4276
rect 8812 4236 9036 4264
rect 8812 4224 8818 4236
rect 9030 4224 9036 4236
rect 9088 4264 9094 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 9088 4236 9137 4264
rect 9088 4224 9094 4236
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9125 4227 9183 4233
rect 10134 4224 10140 4276
rect 10192 4264 10198 4276
rect 13538 4264 13544 4276
rect 10192 4236 13544 4264
rect 10192 4224 10198 4236
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 8312 4196 8340 4224
rect 6932 4168 7696 4196
rect 8312 4168 9352 4196
rect 5276 4126 5856 4128
rect 5215 4100 5856 4126
rect 5215 4098 5304 4100
rect 5215 4097 5227 4098
rect 5169 4091 5227 4097
rect 5902 4088 5908 4140
rect 5960 4088 5966 4140
rect 5997 4132 6055 4137
rect 5997 4131 6224 4132
rect 5997 4097 6009 4131
rect 6043 4128 6224 4131
rect 7006 4128 7012 4140
rect 6043 4104 7012 4128
rect 6043 4097 6055 4104
rect 6196 4100 7012 4104
rect 5997 4091 6055 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7668 4137 7696 4168
rect 7653 4131 7711 4137
rect 7377 4115 7435 4121
rect 7377 4081 7389 4115
rect 7423 4112 7435 4115
rect 7484 4112 7604 4128
rect 7423 4100 7604 4112
rect 7423 4084 7512 4100
rect 7423 4081 7435 4084
rect 7377 4075 7435 4081
rect 6457 4063 6515 4069
rect 5092 4032 5856 4060
rect 4985 4023 5043 4029
rect 3160 3964 4568 3992
rect 1535 3961 1547 3964
rect 1489 3955 1547 3961
rect 1946 3884 1952 3936
rect 2004 3884 2010 3936
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 2556 3896 2605 3924
rect 2556 3884 2562 3896
rect 2593 3893 2605 3896
rect 2639 3924 2651 3927
rect 2866 3924 2872 3936
rect 2639 3896 2872 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 4540 3924 4568 3964
rect 4614 3952 4620 4004
rect 4672 3952 4678 4004
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 5718 3992 5724 4004
rect 4755 3964 5724 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 5828 3992 5856 4032
rect 6457 4029 6469 4063
rect 6503 4060 6515 4063
rect 6546 4060 6552 4072
rect 6503 4032 6552 4060
rect 6503 4029 6515 4032
rect 6457 4023 6515 4029
rect 6546 4020 6552 4032
rect 6604 4060 6610 4072
rect 7098 4060 7104 4072
rect 6604 4032 7104 4060
rect 6604 4020 6610 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7190 4020 7196 4072
rect 7248 4020 7254 4072
rect 7208 3992 7236 4020
rect 5828 3964 7236 3992
rect 7116 3936 7144 3964
rect 4798 3924 4804 3936
rect 4540 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 6089 3927 6147 3933
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 6270 3924 6276 3936
rect 6135 3896 6276 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 7098 3884 7104 3936
rect 7156 3884 7162 3936
rect 7190 3884 7196 3936
rect 7248 3884 7254 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7466 3924 7472 3936
rect 7340 3896 7472 3924
rect 7340 3884 7346 3896
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7576 3924 7604 4100
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 7653 4091 7711 4097
rect 8220 4100 8677 4128
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7800 4032 7849 4060
rect 7800 4020 7806 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8220 3992 8248 4100
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 8478 4020 8484 4072
rect 8536 4020 8542 4072
rect 9324 4060 9352 4168
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 10594 4196 10600 4208
rect 9916 4168 10600 4196
rect 9916 4156 9922 4168
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 11422 4196 11428 4208
rect 10888 4168 11428 4196
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9456 4100 9689 4128
rect 9456 4088 9462 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9944 4131 10002 4137
rect 9944 4097 9956 4131
rect 9990 4128 10002 4131
rect 10888 4128 10916 4168
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 11532 4168 13308 4196
rect 9990 4100 10916 4128
rect 9990 4097 10002 4100
rect 9944 4091 10002 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11296 4100 11345 4128
rect 11296 4088 11302 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11532 4128 11560 4168
rect 11333 4091 11391 4097
rect 11440 4100 11560 4128
rect 12897 4131 12955 4137
rect 11440 4060 11468 4100
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13078 4128 13084 4140
rect 12943 4100 13084 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 9324 4032 9674 4060
rect 7708 3964 8248 3992
rect 7708 3952 7714 3964
rect 8570 3952 8576 4004
rect 8628 3992 8634 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8628 3964 9321 3992
rect 8628 3952 8634 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9030 3924 9036 3936
rect 7576 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9646 3924 9674 4032
rect 10704 4032 11468 4060
rect 10704 3924 10732 4032
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 11974 4060 11980 4072
rect 11756 4032 11980 4060
rect 11756 4020 11762 4032
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 12124 4032 12265 4060
rect 12124 4020 12130 4032
rect 12253 4029 12265 4032
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 11057 3995 11115 4001
rect 11057 3961 11069 3995
rect 11103 3961 11115 3995
rect 11057 3955 11115 3961
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 13188 3992 13216 4091
rect 13280 4069 13308 4168
rect 13998 4156 14004 4208
rect 14056 4196 14062 4208
rect 14093 4199 14151 4205
rect 14093 4196 14105 4199
rect 14056 4168 14105 4196
rect 14056 4156 14062 4168
rect 14093 4165 14105 4168
rect 14139 4165 14151 4199
rect 14093 4159 14151 4165
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13412 4100 13461 4128
rect 13412 4088 13418 4100
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 11195 3964 11468 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 9646 3896 10732 3924
rect 11072 3924 11100 3955
rect 11330 3924 11336 3936
rect 11072 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11440 3924 11468 3964
rect 11624 3964 13216 3992
rect 11624 3924 11652 3964
rect 11440 3896 11652 3924
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11756 3896 12173 3924
rect 11756 3884 11762 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12676 3896 13001 3924
rect 12676 3884 12682 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 14182 3884 14188 3936
rect 14240 3884 14246 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 1118 3680 1124 3732
rect 1176 3720 1182 3732
rect 1765 3723 1823 3729
rect 1765 3720 1777 3723
rect 1176 3692 1777 3720
rect 1176 3680 1182 3692
rect 1765 3689 1777 3692
rect 1811 3689 1823 3723
rect 1765 3683 1823 3689
rect 1854 3680 1860 3732
rect 1912 3680 1918 3732
rect 2498 3680 2504 3732
rect 2556 3680 2562 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3142 3720 3148 3732
rect 2832 3692 3148 3720
rect 2832 3680 2838 3692
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3694 3720 3700 3732
rect 3651 3692 3700 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 4154 3680 4160 3732
rect 4212 3680 4218 3732
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4304 3692 4629 3720
rect 4304 3680 4310 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6638 3720 6644 3732
rect 6319 3692 6644 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7742 3720 7748 3732
rect 7156 3692 7748 3720
rect 7156 3680 7162 3692
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 7892 3692 11376 3720
rect 7892 3680 7898 3692
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 1636 3624 1716 3652
rect 1636 3612 1642 3624
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1688 3516 1716 3624
rect 1872 3584 1900 3680
rect 3786 3652 3792 3664
rect 2148 3624 3792 3652
rect 2041 3587 2099 3593
rect 2041 3584 2053 3587
rect 1872 3556 2053 3584
rect 2041 3553 2053 3556
rect 2087 3553 2099 3587
rect 2041 3547 2099 3553
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1688 3488 1869 3516
rect 1581 3479 1639 3485
rect 1857 3485 1869 3488
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 1596 3448 1624 3479
rect 2148 3448 2176 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 4172 3652 4200 3680
rect 4341 3655 4399 3661
rect 4341 3652 4353 3655
rect 4172 3624 4353 3652
rect 4341 3621 4353 3624
rect 4387 3621 4399 3655
rect 4341 3615 4399 3621
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7524 3624 8156 3652
rect 7524 3612 7530 3624
rect 2976 3593 3280 3596
rect 2959 3587 3280 3593
rect 2959 3553 2971 3587
rect 3005 3584 3280 3587
rect 4065 3587 4123 3593
rect 3005 3568 3924 3584
rect 3005 3553 3017 3568
rect 3252 3556 3924 3568
rect 2959 3547 3017 3553
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2774 3516 2780 3528
rect 2731 3488 2780 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3896 3525 3924 3556
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4246 3584 4252 3596
rect 4111 3556 4252 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4706 3544 4712 3596
rect 4764 3544 4770 3596
rect 8128 3593 8156 3624
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 10594 3652 10600 3664
rect 10468 3624 10600 3652
rect 10468 3612 10474 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 10686 3612 10692 3664
rect 10744 3612 10750 3664
rect 11348 3652 11376 3692
rect 11422 3680 11428 3732
rect 11480 3680 11486 3732
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 11606 3720 11612 3732
rect 11563 3692 11612 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12066 3720 12072 3732
rect 11900 3692 12072 3720
rect 11900 3652 11928 3692
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14148 3692 14289 3720
rect 14148 3680 14154 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 13265 3655 13323 3661
rect 13265 3652 13277 3655
rect 11348 3624 11928 3652
rect 12912 3624 13277 3652
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8202 3584 8208 3596
rect 8159 3556 8208 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 8352 3556 8401 3584
rect 8352 3544 8358 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 11882 3584 11888 3596
rect 10612 3556 10916 3584
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 4724 3516 4752 3544
rect 3927 3488 4752 3516
rect 4801 3519 4859 3525
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 4982 3516 4988 3528
rect 4939 3488 4988 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 3160 3448 3188 3479
rect 1596 3420 2176 3448
rect 2240 3420 3188 3448
rect 750 3340 756 3392
rect 808 3380 814 3392
rect 2240 3380 2268 3420
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4614 3448 4620 3460
rect 3752 3420 4620 3448
rect 3752 3408 3758 3420
rect 4614 3408 4620 3420
rect 4672 3448 4678 3460
rect 4816 3448 4844 3479
rect 4982 3476 4988 3488
rect 5040 3516 5046 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5040 3488 6377 3516
rect 5040 3476 5046 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9398 3516 9404 3528
rect 9355 3488 9404 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9398 3476 9404 3488
rect 9456 3516 9462 3528
rect 10612 3516 10640 3556
rect 9456 3488 10640 3516
rect 9456 3476 9462 3488
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 10744 3488 10793 3516
rect 10744 3476 10750 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10888 3516 10916 3556
rect 11072 3556 11888 3584
rect 11072 3516 11100 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 10888 3488 11100 3516
rect 10781 3479 10839 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11664 3488 11713 3516
rect 11664 3476 11670 3488
rect 11701 3485 11713 3488
rect 11747 3516 11759 3519
rect 12912 3516 12940 3624
rect 13265 3621 13277 3624
rect 13311 3621 13323 3655
rect 13265 3615 13323 3621
rect 14366 3584 14372 3596
rect 11747 3488 12940 3516
rect 13188 3556 14372 3584
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 4672 3420 4844 3448
rect 5160 3451 5218 3457
rect 4672 3408 4678 3420
rect 5160 3417 5172 3451
rect 5206 3448 5218 3451
rect 5810 3448 5816 3460
rect 5206 3420 5816 3448
rect 5206 3417 5218 3420
rect 5160 3411 5218 3417
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 6632 3451 6690 3457
rect 6632 3417 6644 3451
rect 6678 3448 6690 3451
rect 7006 3448 7012 3460
rect 6678 3420 7012 3448
rect 6678 3417 6690 3420
rect 6632 3411 6690 3417
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 8205 3451 8263 3457
rect 7156 3420 7972 3448
rect 7156 3408 7162 3420
rect 808 3352 2268 3380
rect 2777 3383 2835 3389
rect 808 3340 814 3352
rect 2777 3349 2789 3383
rect 2823 3380 2835 3383
rect 7834 3380 7840 3392
rect 2823 3352 7840 3380
rect 2823 3349 2835 3352
rect 2777 3343 2835 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 7944 3380 7972 3420
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 8570 3448 8576 3460
rect 8251 3420 8576 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 9576 3451 9634 3457
rect 9576 3417 9588 3451
rect 9622 3448 9634 3451
rect 11882 3448 11888 3460
rect 9622 3420 11888 3448
rect 9622 3417 9634 3420
rect 9576 3411 9634 3417
rect 11882 3408 11888 3420
rect 11940 3408 11946 3460
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 12130 3451 12188 3457
rect 12130 3448 12142 3451
rect 12032 3420 12142 3448
rect 12032 3408 12038 3420
rect 12130 3417 12142 3420
rect 12176 3417 12188 3451
rect 13188 3448 13216 3556
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 13446 3476 13452 3528
rect 13504 3476 13510 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13780 3488 14105 3516
rect 13780 3476 13786 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 12130 3411 12188 3417
rect 12406 3420 13216 3448
rect 13817 3451 13875 3457
rect 12406 3380 12434 3420
rect 13817 3417 13829 3451
rect 13863 3448 13875 3451
rect 14550 3448 14556 3460
rect 13863 3420 14556 3448
rect 13863 3417 13875 3420
rect 13817 3411 13875 3417
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 7944 3352 12434 3380
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 2314 3176 2320 3188
rect 2179 3148 2320 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3326 3176 3332 3188
rect 3283 3148 3332 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 4062 3176 4068 3188
rect 3467 3148 4068 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 4212 3148 4261 3176
rect 4212 3136 4218 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 5074 3176 5080 3188
rect 4479 3148 5080 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6546 3136 6552 3188
rect 6604 3136 6610 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7248 3148 8892 3176
rect 7248 3136 7254 3148
rect 3878 3068 3884 3120
rect 3936 3108 3942 3120
rect 6564 3108 6592 3136
rect 3936 3080 4384 3108
rect 6564 3080 6868 3108
rect 3936 3068 3942 3080
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1360 3012 1409 3040
rect 1360 3000 1366 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2777 3043 2835 3049
rect 2271 3012 2728 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 474 2932 480 2984
rect 532 2932 538 2984
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 1964 2972 1992 3003
rect 624 2944 1992 2972
rect 624 2932 630 2944
rect 492 2836 520 2932
rect 1486 2864 1492 2916
rect 1544 2864 1550 2916
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 492 2808 1869 2836
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 1857 2799 1915 2805
rect 2406 2796 2412 2848
rect 2464 2796 2470 2848
rect 2700 2836 2728 3012
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2823 3012 3065 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3068 2972 3096 3003
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3292 3012 3341 3040
rect 3292 3000 3298 3012
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3568 3012 3617 3040
rect 3568 3000 3574 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 4062 3040 4068 3052
rect 3605 3003 3663 3009
rect 3712 3012 4068 3040
rect 3712 2972 3740 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4356 3049 4384 3080
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4798 3000 4804 3052
rect 4856 3000 4862 3052
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3040 6515 3043
rect 6638 3040 6644 3052
rect 6503 3012 6644 3040
rect 6503 3009 6515 3012
rect 6457 3003 6515 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6730 3000 6736 3052
rect 6788 3000 6794 3052
rect 3068 2944 3740 2972
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 3804 2904 3832 2935
rect 5534 2932 5540 2984
rect 5592 2932 5598 2984
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6748 2972 6776 3000
rect 5767 2944 6776 2972
rect 6840 2972 6868 3080
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 7285 3111 7343 3117
rect 7285 3108 7297 3111
rect 6972 3080 7297 3108
rect 6972 3068 6978 3080
rect 7285 3077 7297 3080
rect 7331 3077 7343 3111
rect 7285 3071 7343 3077
rect 7650 3068 7656 3120
rect 7708 3108 7714 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7708 3080 7849 3108
rect 7708 3068 7714 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 8573 3111 8631 3117
rect 8573 3108 8585 3111
rect 8260 3080 8585 3108
rect 8260 3068 8266 3080
rect 8573 3077 8585 3080
rect 8619 3077 8631 3111
rect 8573 3071 8631 3077
rect 8754 3068 8760 3120
rect 8812 3068 8818 3120
rect 8864 3117 8892 3148
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9088 3148 9505 3176
rect 9088 3136 9094 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 11238 3176 11244 3188
rect 9640 3148 11244 3176
rect 9640 3136 9646 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11698 3136 11704 3188
rect 11756 3136 11762 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11940 3148 12173 3176
rect 11940 3136 11946 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 12308 3148 12388 3176
rect 12308 3136 12314 3148
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3077 8907 3111
rect 8849 3071 8907 3077
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 10128 3111 10186 3117
rect 9272 3080 9720 3108
rect 9272 3068 9278 3080
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 9692 3049 9720 3080
rect 10128 3077 10140 3111
rect 10174 3108 10186 3111
rect 11716 3108 11744 3136
rect 12360 3117 12388 3148
rect 13630 3136 13636 3188
rect 13688 3136 13694 3188
rect 10174 3080 10824 3108
rect 10174 3077 10186 3080
rect 10128 3071 10186 3077
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 10686 3040 10692 3052
rect 9677 3003 9735 3009
rect 9784 3012 10692 3040
rect 6840 2944 7144 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 3016 2876 3832 2904
rect 3016 2864 3022 2876
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 6181 2907 6239 2913
rect 4028 2876 6132 2904
rect 4028 2864 4034 2876
rect 4338 2836 4344 2848
rect 2700 2808 4344 2836
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5534 2836 5540 2848
rect 5491 2808 5540 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6104 2836 6132 2876
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 7006 2904 7012 2916
rect 6227 2876 7012 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7116 2904 7144 2944
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7374 2972 7380 2984
rect 7248 2944 7380 2972
rect 7248 2932 7254 2944
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8110 2932 8116 2984
rect 8168 2932 8174 2984
rect 8312 2972 8340 3000
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8312 2944 9045 2972
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9582 2972 9588 2984
rect 9033 2935 9091 2941
rect 9140 2944 9588 2972
rect 9140 2904 9168 2944
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 7116 2876 9168 2904
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 9784 2904 9812 3012
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10796 3040 10824 3080
rect 11164 3080 11744 3108
rect 12345 3111 12403 3117
rect 11164 3040 11192 3080
rect 12345 3077 12357 3111
rect 12391 3077 12403 3111
rect 12345 3071 12403 3077
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3108 12495 3111
rect 12526 3108 12532 3120
rect 12483 3080 12532 3108
rect 12483 3077 12495 3080
rect 12437 3071 12495 3077
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 12989 3111 13047 3117
rect 12989 3077 13001 3111
rect 13035 3108 13047 3111
rect 13354 3108 13360 3120
rect 13035 3080 13360 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 13354 3068 13360 3080
rect 13412 3108 13418 3120
rect 13648 3108 13676 3136
rect 13412 3080 13676 3108
rect 13412 3068 13418 3080
rect 10796 3012 11192 3040
rect 11606 3000 11612 3052
rect 11664 3000 11670 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 14458 3040 14464 3052
rect 13679 3012 14464 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 9272 2876 9812 2904
rect 9272 2864 9278 2876
rect 7926 2836 7932 2848
rect 6104 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9876 2836 9904 2935
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 12158 2972 12164 2984
rect 10928 2944 12164 2972
rect 10928 2932 10934 2944
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13188 2972 13216 3003
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 12768 2944 13216 2972
rect 13909 2975 13967 2981
rect 12768 2932 12774 2944
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 14366 2972 14372 2984
rect 13955 2944 14372 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 11606 2864 11612 2916
rect 11664 2904 11670 2916
rect 13814 2904 13820 2916
rect 11664 2876 13820 2904
rect 11664 2864 11670 2876
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 9456 2808 9904 2836
rect 9456 2796 9462 2808
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 10192 2808 13277 2836
rect 10192 2796 10198 2808
rect 13265 2805 13277 2808
rect 13311 2805 13323 2839
rect 13265 2799 13323 2805
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 382 2592 388 2644
rect 440 2632 446 2644
rect 2498 2632 2504 2644
rect 440 2604 2504 2632
rect 440 2592 446 2604
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3050 2632 3056 2644
rect 2823 2604 3056 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 4433 2635 4491 2641
rect 3528 2604 3740 2632
rect 658 2524 664 2576
rect 716 2564 722 2576
rect 2409 2567 2467 2573
rect 716 2536 2176 2564
rect 716 2524 722 2536
rect 1394 2456 1400 2508
rect 1452 2456 1458 2508
rect 2148 2496 2176 2536
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 3528 2564 3556 2604
rect 2455 2536 3556 2564
rect 3605 2567 3663 2573
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 3605 2533 3617 2567
rect 3651 2533 3663 2567
rect 3605 2527 3663 2533
rect 3620 2496 3648 2527
rect 2148 2468 3648 2496
rect 3712 2496 3740 2604
rect 4172 2604 4384 2632
rect 4172 2573 4200 2604
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2533 4215 2567
rect 4356 2564 4384 2604
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 5074 2632 5080 2644
rect 4479 2604 5080 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 9674 2632 9680 2644
rect 7892 2604 9680 2632
rect 7892 2592 7898 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10502 2632 10508 2644
rect 9815 2604 10508 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 12802 2632 12808 2644
rect 11379 2604 12808 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 14093 2635 14151 2641
rect 12912 2604 13860 2632
rect 4798 2564 4804 2576
rect 4356 2536 4804 2564
rect 4157 2527 4215 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 4985 2567 5043 2573
rect 4985 2533 4997 2567
rect 5031 2564 5043 2567
rect 5031 2536 8432 2564
rect 5031 2533 5043 2536
rect 4985 2527 5043 2533
rect 5169 2499 5227 2505
rect 3712 2468 4292 2496
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2280 2400 2329 2428
rect 2280 2388 2286 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 2884 2360 2912 2391
rect 3142 2388 3148 2440
rect 3200 2388 3206 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 3292 2400 3433 2428
rect 3292 2388 3298 2400
rect 3421 2397 3433 2400
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 3694 2360 3700 2372
rect 2884 2332 3700 2360
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 2958 2252 2964 2304
rect 3016 2252 3022 2304
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 3970 2252 3976 2304
rect 4028 2252 4034 2304
rect 4080 2292 4108 2391
rect 4264 2360 4292 2468
rect 4540 2468 5028 2496
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4540 2428 4568 2468
rect 4396 2400 4568 2428
rect 4396 2388 4402 2400
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 5000 2428 5028 2468
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5442 2496 5448 2508
rect 5215 2468 5448 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 5592 2468 7021 2496
rect 5592 2456 5598 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7650 2456 7656 2508
rect 7708 2456 7714 2508
rect 8110 2456 8116 2508
rect 8168 2456 8174 2508
rect 5258 2428 5264 2440
rect 5000 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 6454 2388 6460 2440
rect 6512 2388 6518 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 5644 2360 5672 2388
rect 4264 2332 5672 2360
rect 5997 2363 6055 2369
rect 5997 2329 6009 2363
rect 6043 2360 6055 2363
rect 6043 2332 7052 2360
rect 6043 2329 6055 2332
rect 5997 2323 6055 2329
rect 4522 2292 4528 2304
rect 4080 2264 4528 2292
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 6638 2292 6644 2304
rect 5316 2264 6644 2292
rect 5316 2252 5322 2264
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 6730 2252 6736 2304
rect 6788 2252 6794 2304
rect 7024 2292 7052 2332
rect 7098 2320 7104 2372
rect 7156 2320 7162 2372
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 8128 2360 8156 2456
rect 8404 2437 8432 2536
rect 8570 2524 8576 2576
rect 8628 2564 8634 2576
rect 10597 2567 10655 2573
rect 8628 2536 9996 2564
rect 8628 2524 8634 2536
rect 9766 2496 9772 2508
rect 8496 2468 9772 2496
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 7248 2332 8156 2360
rect 8220 2360 8248 2391
rect 8496 2360 8524 2468
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9723 2400 9904 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 8220 2332 8524 2360
rect 7248 2320 7254 2332
rect 8570 2320 8576 2372
rect 8628 2320 8634 2372
rect 8757 2363 8815 2369
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 9398 2360 9404 2372
rect 8803 2332 9404 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 8588 2292 8616 2320
rect 7024 2264 8616 2292
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8720 2264 9137 2292
rect 8720 2252 8726 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9876 2292 9904 2400
rect 9968 2360 9996 2536
rect 10597 2533 10609 2567
rect 10643 2564 10655 2567
rect 11974 2564 11980 2576
rect 10643 2536 11980 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 12912 2564 12940 2604
rect 12406 2536 12940 2564
rect 12989 2567 13047 2573
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10376 2468 10701 2496
rect 10376 2456 10382 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 10778 2456 10784 2508
rect 10836 2496 10842 2508
rect 10873 2499 10931 2505
rect 10873 2496 10885 2499
rect 10836 2468 10885 2496
rect 10836 2456 10842 2468
rect 10873 2465 10885 2468
rect 10919 2465 10931 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 10873 2459 10931 2465
rect 11164 2468 11897 2496
rect 11164 2440 11192 2468
rect 11885 2465 11897 2468
rect 11931 2496 11943 2499
rect 12406 2496 12434 2536
rect 12989 2533 13001 2567
rect 13035 2564 13047 2567
rect 13354 2564 13360 2576
rect 13035 2536 13360 2564
rect 13035 2533 13047 2536
rect 12989 2527 13047 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 13832 2573 13860 2604
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14274 2632 14280 2644
rect 14139 2604 14280 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 13817 2567 13875 2573
rect 13817 2533 13829 2567
rect 13863 2533 13875 2567
rect 13817 2527 13875 2533
rect 11931 2468 12434 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 13262 2496 13268 2508
rect 12860 2468 13268 2496
rect 12860 2456 12866 2468
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10410 2428 10416 2440
rect 10091 2424 10171 2428
rect 10244 2424 10416 2428
rect 10091 2400 10416 2424
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10143 2396 10272 2400
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 14274 2388 14280 2440
rect 14332 2388 14338 2440
rect 11609 2363 11667 2369
rect 11609 2360 11621 2363
rect 9968 2332 11621 2360
rect 11609 2329 11621 2332
rect 11655 2329 11667 2363
rect 11609 2323 11667 2329
rect 11698 2320 11704 2372
rect 11756 2320 11762 2372
rect 11882 2320 11888 2372
rect 11940 2320 11946 2372
rect 12434 2320 12440 2372
rect 12492 2320 12498 2372
rect 12526 2320 12532 2372
rect 12584 2320 12590 2372
rect 13357 2363 13415 2369
rect 13357 2329 13369 2363
rect 13403 2329 13415 2363
rect 13357 2323 13415 2329
rect 10962 2292 10968 2304
rect 9876 2264 10968 2292
rect 9125 2255 9183 2261
rect 10962 2252 10968 2264
rect 11020 2292 11026 2304
rect 11900 2292 11928 2320
rect 11020 2264 11928 2292
rect 11020 2252 11026 2264
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 13372 2292 13400 2323
rect 12216 2264 13400 2292
rect 12216 2252 12222 2264
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 1670 2048 1676 2100
rect 1728 2048 1734 2100
rect 2406 2048 2412 2100
rect 2464 2048 2470 2100
rect 3786 2088 3792 2100
rect 2746 2060 3792 2088
rect 1688 1816 1716 2048
rect 2424 2020 2452 2048
rect 2746 2020 2774 2060
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 13078 2088 13084 2100
rect 6788 2060 13084 2088
rect 6788 2048 6794 2060
rect 13078 2048 13084 2060
rect 13136 2048 13142 2100
rect 2424 1992 2774 2020
rect 4890 1980 4896 2032
rect 4948 2020 4954 2032
rect 8294 2020 8300 2032
rect 4948 1992 8300 2020
rect 4948 1980 4954 1992
rect 8294 1980 8300 1992
rect 8352 1980 8358 2032
rect 8478 1980 8484 2032
rect 8536 1980 8542 2032
rect 8754 1980 8760 2032
rect 8812 1980 8818 2032
rect 9950 1980 9956 2032
rect 10008 2020 10014 2032
rect 12158 2020 12164 2032
rect 10008 1992 12164 2020
rect 10008 1980 10014 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 4706 1912 4712 1964
rect 4764 1952 4770 1964
rect 8496 1952 8524 1980
rect 4764 1924 8524 1952
rect 8772 1952 8800 1980
rect 11146 1952 11152 1964
rect 8772 1924 11152 1952
rect 4764 1912 4770 1924
rect 11146 1912 11152 1924
rect 11204 1912 11210 1964
rect 4798 1844 4804 1896
rect 4856 1884 4862 1896
rect 12710 1884 12716 1896
rect 4856 1856 12716 1884
rect 4856 1844 4862 1856
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 1688 1788 2774 1816
rect 2746 1748 2774 1788
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 7190 1816 7196 1828
rect 3016 1788 7196 1816
rect 3016 1776 3022 1788
rect 7190 1776 7196 1788
rect 7248 1776 7254 1828
rect 9766 1816 9772 1828
rect 7300 1788 9772 1816
rect 2746 1720 3004 1748
rect 2976 1680 3004 1720
rect 3970 1708 3976 1760
rect 4028 1748 4034 1760
rect 7300 1748 7328 1788
rect 9766 1776 9772 1788
rect 9824 1776 9830 1828
rect 4028 1720 7328 1748
rect 4028 1708 4034 1720
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 11238 1748 11244 1760
rect 8260 1720 11244 1748
rect 8260 1708 8266 1720
rect 11238 1708 11244 1720
rect 11296 1708 11302 1760
rect 8938 1680 8944 1692
rect 2976 1652 8944 1680
rect 8938 1640 8944 1652
rect 8996 1640 9002 1692
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 9950 1340 9956 1352
rect 5040 1312 9956 1340
rect 5040 1300 5046 1312
rect 9950 1300 9956 1312
rect 10008 1300 10014 1352
rect 10226 1232 10232 1284
rect 10284 1272 10290 1284
rect 12342 1272 12348 1284
rect 10284 1244 12348 1272
rect 10284 1232 10290 1244
rect 12342 1232 12348 1244
rect 12400 1232 12406 1284
<< via1 >>
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 13728 17280 13780 17332
rect 14556 17280 14608 17332
rect 2780 17255 2832 17264
rect 2780 17221 2789 17255
rect 2789 17221 2823 17255
rect 2823 17221 2832 17255
rect 2780 17212 2832 17221
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 10968 17144 11020 17196
rect 5632 17076 5684 17128
rect 1032 16940 1084 16992
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 940 16736 992 16788
rect 2412 16736 2464 16788
rect 14648 16736 14700 16788
rect 9864 16600 9916 16652
rect 8760 16532 8812 16584
rect 15016 16532 15068 16584
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 13820 16396 13872 16448
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 940 16192 992 16244
rect 9956 16056 10008 16108
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 1124 15648 1176 15700
rect 3424 15444 3476 15496
rect 13820 15648 13872 15700
rect 14832 15580 14884 15632
rect 13912 15444 13964 15496
rect 2872 15376 2924 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 5908 15308 5960 15360
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 1676 14968 1728 15020
rect 8208 15104 8260 15156
rect 7196 15036 7248 15088
rect 9956 15036 10008 15088
rect 12072 15036 12124 15088
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 4896 14968 4948 15020
rect 10784 14968 10836 15020
rect 4160 14900 4212 14952
rect 3608 14832 3660 14884
rect 1400 14807 1452 14816
rect 1400 14773 1409 14807
rect 1409 14773 1443 14807
rect 1443 14773 1452 14807
rect 1400 14764 1452 14773
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 3240 14807 3292 14816
rect 3240 14773 3249 14807
rect 3249 14773 3283 14807
rect 3283 14773 3292 14807
rect 3240 14764 3292 14773
rect 3332 14764 3384 14816
rect 9128 14764 9180 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 1400 14560 1452 14612
rect 1860 14356 1912 14408
rect 2412 14467 2464 14476
rect 2412 14433 2421 14467
rect 2421 14433 2455 14467
rect 2455 14433 2464 14467
rect 2412 14424 2464 14433
rect 3516 14560 3568 14612
rect 10232 14560 10284 14612
rect 9864 14492 9916 14544
rect 2964 14356 3016 14408
rect 3700 14424 3752 14476
rect 9956 14424 10008 14476
rect 3516 14356 3568 14408
rect 8300 14356 8352 14408
rect 3792 14288 3844 14340
rect 9312 14288 9364 14340
rect 9496 14331 9548 14340
rect 9496 14297 9505 14331
rect 9505 14297 9539 14331
rect 9539 14297 9548 14331
rect 9496 14288 9548 14297
rect 1860 14220 1912 14272
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 3516 14220 3568 14272
rect 5264 14220 5316 14272
rect 8392 14263 8444 14272
rect 8392 14229 8401 14263
rect 8401 14229 8435 14263
rect 8435 14229 8444 14263
rect 8392 14220 8444 14229
rect 8484 14220 8536 14272
rect 10968 14356 11020 14408
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 1216 14016 1268 14068
rect 3056 14016 3108 14068
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 1492 13991 1544 14000
rect 1492 13957 1501 13991
rect 1501 13957 1535 13991
rect 1535 13957 1544 13991
rect 1492 13948 1544 13957
rect 1676 13948 1728 14000
rect 480 13880 532 13932
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 2504 13880 2556 13932
rect 3700 14016 3752 14068
rect 5080 14016 5132 14068
rect 8576 14059 8628 14068
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 9496 14016 9548 14068
rect 10968 14016 11020 14068
rect 13728 14016 13780 14068
rect 3792 13948 3844 14000
rect 4804 13948 4856 14000
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 756 13744 808 13796
rect 3424 13744 3476 13796
rect 3516 13744 3568 13796
rect 3792 13812 3844 13864
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 6920 13812 6972 13864
rect 7656 13812 7708 13864
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 9220 13812 9272 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 14464 13812 14516 13864
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 3240 13676 3292 13728
rect 3332 13676 3384 13728
rect 10876 13744 10928 13796
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 12716 13719 12768 13728
rect 12716 13685 12725 13719
rect 12725 13685 12759 13719
rect 12759 13685 12768 13719
rect 12716 13676 12768 13685
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 1124 13404 1176 13456
rect 572 13336 624 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 3240 13336 3292 13388
rect 664 13200 716 13252
rect 3332 13268 3384 13320
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 2964 13200 3016 13252
rect 940 13132 992 13184
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 3608 13175 3660 13184
rect 3608 13141 3617 13175
rect 3617 13141 3651 13175
rect 3651 13141 3660 13175
rect 3608 13132 3660 13141
rect 6000 13200 6052 13252
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 8116 13472 8168 13524
rect 8300 13472 8352 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 8760 13472 8812 13524
rect 10324 13515 10376 13524
rect 10324 13481 10333 13515
rect 10333 13481 10367 13515
rect 10367 13481 10376 13515
rect 10324 13472 10376 13481
rect 14280 13472 14332 13524
rect 8392 13336 8444 13388
rect 8484 13268 8536 13320
rect 11060 13268 11112 13320
rect 12716 13336 12768 13388
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 8392 13200 8444 13252
rect 8668 13200 8720 13252
rect 9312 13200 9364 13252
rect 12256 13200 12308 13252
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 11612 13132 11664 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 2136 12928 2188 12980
rect 388 12860 440 12912
rect 4252 12860 4304 12912
rect 4528 12860 4580 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 2044 12792 2096 12844
rect 2964 12792 3016 12844
rect 848 12588 900 12640
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2412 12588 2464 12640
rect 2964 12656 3016 12708
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 7104 12860 7156 12912
rect 8576 12928 8628 12980
rect 11796 12928 11848 12980
rect 12992 12928 13044 12980
rect 4068 12724 4120 12776
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4344 12724 4396 12776
rect 5264 12724 5316 12776
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 7288 12792 7340 12844
rect 5816 12767 5868 12776
rect 5816 12733 5825 12767
rect 5825 12733 5859 12767
rect 5859 12733 5868 12767
rect 5816 12724 5868 12733
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 8300 12724 8352 12776
rect 3240 12588 3292 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 6644 12588 6696 12640
rect 8392 12656 8444 12708
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 10416 12792 10468 12844
rect 11520 12860 11572 12912
rect 12624 12860 12676 12912
rect 9036 12656 9088 12708
rect 8668 12588 8720 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 12716 12656 12768 12708
rect 12440 12588 12492 12640
rect 13268 12588 13320 12640
rect 13544 12588 13596 12640
rect 14464 12724 14516 12776
rect 14556 12588 14608 12640
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 2504 12384 2556 12436
rect 3424 12384 3476 12436
rect 4068 12384 4120 12436
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 3516 12248 3568 12300
rect 3884 12248 3936 12300
rect 4160 12316 4212 12368
rect 4344 12248 4396 12300
rect 1492 12155 1544 12164
rect 1492 12121 1501 12155
rect 1501 12121 1535 12155
rect 1535 12121 1544 12155
rect 1492 12112 1544 12121
rect 2504 12112 2556 12164
rect 2872 12112 2924 12164
rect 940 12044 992 12096
rect 3240 12044 3292 12096
rect 3424 12044 3476 12096
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 5540 12180 5592 12232
rect 6736 12248 6788 12300
rect 7196 12248 7248 12300
rect 9220 12384 9272 12436
rect 12992 12384 13044 12436
rect 13452 12384 13504 12436
rect 14188 12384 14240 12436
rect 6000 12180 6052 12232
rect 6828 12180 6880 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 12164 12291 12216 12300
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 12164 12248 12216 12257
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 14372 12359 14424 12368
rect 14372 12325 14381 12359
rect 14381 12325 14415 12359
rect 14415 12325 14424 12359
rect 14372 12316 14424 12325
rect 4160 12155 4212 12164
rect 4160 12121 4169 12155
rect 4169 12121 4203 12155
rect 4203 12121 4212 12155
rect 4160 12112 4212 12121
rect 4528 12112 4580 12164
rect 5356 12112 5408 12164
rect 4712 12044 4764 12096
rect 5632 12044 5684 12096
rect 8484 12180 8536 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9036 12180 9088 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 11152 12180 11204 12232
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 11612 12112 11664 12164
rect 12348 12112 12400 12164
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 10048 12044 10100 12096
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 1492 11840 1544 11892
rect 2872 11840 2924 11892
rect 1676 11704 1728 11756
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2412 11636 2464 11688
rect 1216 11568 1268 11620
rect 1400 11500 1452 11552
rect 1676 11500 1728 11552
rect 2136 11500 2188 11552
rect 3424 11772 3476 11824
rect 3792 11840 3844 11892
rect 3148 11747 3200 11756
rect 3148 11713 3182 11747
rect 3182 11713 3200 11747
rect 3148 11704 3200 11713
rect 4252 11840 4304 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 7564 11840 7616 11892
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 8484 11840 8536 11892
rect 10232 11840 10284 11892
rect 10968 11840 11020 11892
rect 11152 11840 11204 11892
rect 6828 11772 6880 11824
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 6000 11704 6052 11756
rect 7656 11772 7708 11824
rect 8392 11772 8444 11824
rect 7472 11704 7524 11756
rect 10416 11772 10468 11824
rect 2504 11500 2556 11552
rect 4712 11568 4764 11620
rect 5172 11636 5224 11688
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 6920 11636 6972 11688
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 13176 11840 13228 11892
rect 13636 11883 13688 11892
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 14188 11840 14240 11892
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 13268 11704 13320 11756
rect 3976 11500 4028 11552
rect 5724 11500 5776 11552
rect 6828 11611 6880 11620
rect 6828 11577 6837 11611
rect 6837 11577 6871 11611
rect 6871 11577 6880 11611
rect 6828 11568 6880 11577
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 7288 11500 7340 11552
rect 7748 11500 7800 11552
rect 9220 11500 9272 11552
rect 12716 11568 12768 11620
rect 14280 11500 14332 11552
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 1492 11296 1544 11348
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2044 11092 2096 11144
rect 3148 11296 3200 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4068 11296 4120 11348
rect 7380 11296 7432 11348
rect 7472 11296 7524 11348
rect 3608 11228 3660 11280
rect 5724 11228 5776 11280
rect 6552 11228 6604 11280
rect 7288 11228 7340 11280
rect 2780 11092 2832 11144
rect 4068 11092 4120 11144
rect 5540 11092 5592 11144
rect 4252 11024 4304 11076
rect 4804 11024 4856 11076
rect 7748 11228 7800 11280
rect 8944 11296 8996 11348
rect 9220 11228 9272 11280
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 13268 11296 13320 11348
rect 13636 11296 13688 11348
rect 11888 11160 11940 11212
rect 6828 11024 6880 11076
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 8484 11092 8536 11144
rect 8852 11092 8904 11144
rect 11060 11092 11112 11144
rect 12164 11092 12216 11144
rect 13728 11228 13780 11280
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 3056 10956 3108 11008
rect 3148 10956 3200 11008
rect 3608 10956 3660 11008
rect 3976 10956 4028 11008
rect 5540 10956 5592 11008
rect 10416 11024 10468 11076
rect 13360 11024 13412 11076
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 9956 10956 10008 11008
rect 10692 10956 10744 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 13636 10956 13688 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 3332 10752 3384 10804
rect 4068 10752 4120 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 6000 10752 6052 10804
rect 7104 10752 7156 10804
rect 8852 10752 8904 10804
rect 8944 10752 8996 10804
rect 9404 10752 9456 10804
rect 12164 10752 12216 10804
rect 940 10616 992 10668
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 1676 10548 1728 10600
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3240 10616 3292 10668
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 6552 10727 6604 10736
rect 6552 10693 6561 10727
rect 6561 10693 6595 10727
rect 6595 10693 6604 10727
rect 6552 10684 6604 10693
rect 7656 10684 7708 10736
rect 8760 10684 8812 10736
rect 3332 10548 3384 10600
rect 6460 10591 6512 10600
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3976 10412 4028 10464
rect 5540 10412 5592 10464
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 7288 10548 7340 10600
rect 6000 10480 6052 10532
rect 7104 10480 7156 10532
rect 8484 10616 8536 10668
rect 9220 10548 9272 10600
rect 10048 10616 10100 10668
rect 10508 10616 10560 10668
rect 6736 10412 6788 10464
rect 9404 10412 9456 10464
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11060 10616 11112 10668
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 12624 10684 12676 10736
rect 13176 10684 13228 10736
rect 11152 10548 11204 10600
rect 13452 10548 13504 10600
rect 9956 10412 10008 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 12716 10412 12768 10464
rect 13636 10480 13688 10532
rect 14096 10412 14148 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 3792 10208 3844 10260
rect 3976 10208 4028 10260
rect 6000 10208 6052 10260
rect 6184 10208 6236 10260
rect 3424 10140 3476 10192
rect 4896 10140 4948 10192
rect 6368 10140 6420 10192
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 6092 10072 6144 10124
rect 6552 10208 6604 10260
rect 7288 10208 7340 10260
rect 9404 10208 9456 10260
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3700 10004 3752 10056
rect 3884 10004 3936 10056
rect 4252 10004 4304 10056
rect 2136 9936 2188 9988
rect 5724 10004 5776 10056
rect 6920 10072 6972 10124
rect 9220 10115 9272 10124
rect 9220 10081 9229 10115
rect 9229 10081 9263 10115
rect 9263 10081 9272 10115
rect 10048 10208 10100 10260
rect 10876 10208 10928 10260
rect 11336 10208 11388 10260
rect 9220 10072 9272 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10600 10140 10652 10192
rect 5540 9936 5592 9988
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 9312 10004 9364 10056
rect 9680 10004 9732 10056
rect 9772 9936 9824 9988
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 3608 9868 3660 9920
rect 5356 9868 5408 9920
rect 6000 9868 6052 9920
rect 6736 9868 6788 9920
rect 9404 9868 9456 9920
rect 10416 10072 10468 10124
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 13452 10183 13504 10192
rect 13452 10149 13461 10183
rect 13461 10149 13495 10183
rect 13495 10149 13504 10183
rect 13452 10140 13504 10149
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12808 10072 12860 10124
rect 13728 10072 13780 10124
rect 11980 10004 12032 10056
rect 12164 10004 12216 10056
rect 12716 9936 12768 9988
rect 12900 9936 12952 9988
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13176 10004 13228 10056
rect 14464 10004 14516 10056
rect 10968 9868 11020 9920
rect 12164 9868 12216 9920
rect 12624 9868 12676 9920
rect 13636 9868 13688 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 1400 9664 1452 9716
rect 1676 9664 1728 9716
rect 1952 9664 2004 9716
rect 3148 9664 3200 9716
rect 3700 9664 3752 9716
rect 3884 9664 3936 9716
rect 4252 9664 4304 9716
rect 5172 9664 5224 9716
rect 6184 9664 6236 9716
rect 6460 9664 6512 9716
rect 6552 9664 6604 9716
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 3056 9528 3108 9580
rect 3424 9528 3476 9580
rect 6736 9596 6788 9648
rect 1676 9460 1728 9512
rect 1768 9324 1820 9376
rect 3148 9460 3200 9512
rect 6000 9528 6052 9580
rect 6368 9528 6420 9580
rect 5908 9460 5960 9512
rect 5080 9324 5132 9376
rect 5908 9324 5960 9376
rect 6552 9324 6604 9376
rect 6736 9460 6788 9512
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 6920 9392 6972 9444
rect 7104 9596 7156 9648
rect 9404 9664 9456 9716
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 9036 9596 9088 9648
rect 10508 9596 10560 9648
rect 12900 9664 12952 9716
rect 13084 9664 13136 9716
rect 14188 9707 14240 9716
rect 14188 9673 14197 9707
rect 14197 9673 14231 9707
rect 14231 9673 14240 9707
rect 14188 9664 14240 9673
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8300 9460 8352 9512
rect 9128 9460 9180 9512
rect 7656 9392 7708 9444
rect 8576 9435 8628 9444
rect 8576 9401 8585 9435
rect 8585 9401 8619 9435
rect 8619 9401 8628 9435
rect 8576 9392 8628 9401
rect 9312 9392 9364 9444
rect 9496 9435 9548 9444
rect 9496 9401 9505 9435
rect 9505 9401 9539 9435
rect 9539 9401 9548 9435
rect 9496 9392 9548 9401
rect 7932 9367 7984 9376
rect 7932 9333 7941 9367
rect 7941 9333 7975 9367
rect 7975 9333 7984 9367
rect 7932 9324 7984 9333
rect 8668 9324 8720 9376
rect 9772 9528 9824 9580
rect 9772 9392 9824 9444
rect 10048 9324 10100 9376
rect 10416 9528 10468 9580
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 12716 9596 12768 9648
rect 11244 9528 11296 9580
rect 11704 9460 11756 9512
rect 12164 9460 12216 9512
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12808 9528 12860 9580
rect 13360 9639 13412 9648
rect 13360 9605 13369 9639
rect 13369 9605 13403 9639
rect 13403 9605 13412 9639
rect 13360 9596 13412 9605
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 10416 9392 10468 9444
rect 10508 9324 10560 9376
rect 11888 9324 11940 9376
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 11980 9324 12032 9333
rect 13360 9324 13412 9376
rect 13820 9324 13872 9376
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 2412 9120 2464 9172
rect 2688 9120 2740 9172
rect 3148 9120 3200 9172
rect 3976 9120 4028 9172
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 3424 9052 3476 9104
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 940 8916 992 8968
rect 2228 8916 2280 8968
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 6000 9052 6052 9104
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 7656 9120 7708 9172
rect 8300 9120 8352 9172
rect 940 8780 992 8832
rect 1400 8823 1452 8832
rect 1400 8789 1409 8823
rect 1409 8789 1443 8823
rect 1443 8789 1452 8823
rect 1400 8780 1452 8789
rect 2320 8780 2372 8832
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 3148 8848 3200 8900
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 10048 9052 10100 9104
rect 11704 9120 11756 9172
rect 12624 9120 12676 9172
rect 6920 8984 6972 9036
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 10968 9052 11020 9104
rect 11152 8984 11204 9036
rect 14096 9052 14148 9104
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 13360 8984 13412 9036
rect 5172 8848 5224 8900
rect 4252 8780 4304 8832
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6552 8848 6604 8900
rect 6828 8848 6880 8900
rect 6368 8780 6420 8832
rect 7288 8916 7340 8968
rect 8668 8848 8720 8900
rect 7748 8780 7800 8832
rect 9404 8848 9456 8900
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 9772 8780 9824 8832
rect 10508 8780 10560 8832
rect 11060 8780 11112 8832
rect 11888 8916 11940 8968
rect 12900 8916 12952 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 12624 8823 12676 8832
rect 12624 8789 12633 8823
rect 12633 8789 12667 8823
rect 12667 8789 12676 8823
rect 12624 8780 12676 8789
rect 12808 8780 12860 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13544 8780 13596 8832
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 2136 8576 2188 8628
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 3608 8508 3660 8560
rect 2688 8440 2740 8492
rect 3792 8440 3844 8492
rect 4620 8440 4672 8492
rect 4988 8576 5040 8628
rect 6276 8576 6328 8628
rect 6736 8576 6788 8628
rect 7196 8576 7248 8628
rect 9956 8576 10008 8628
rect 5356 8508 5408 8560
rect 6460 8508 6512 8560
rect 1676 8372 1728 8424
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2504 8372 2556 8424
rect 3056 8372 3108 8424
rect 1768 8304 1820 8356
rect 3884 8304 3936 8356
rect 3976 8304 4028 8356
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6736 8440 6788 8492
rect 7380 8551 7432 8560
rect 7380 8517 7389 8551
rect 7389 8517 7423 8551
rect 7423 8517 7432 8551
rect 7380 8508 7432 8517
rect 10324 8576 10376 8628
rect 10416 8576 10468 8628
rect 10784 8576 10836 8628
rect 11704 8576 11756 8628
rect 11888 8576 11940 8628
rect 12624 8576 12676 8628
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 10508 8508 10560 8560
rect 14372 8508 14424 8560
rect 6460 8372 6512 8424
rect 8300 8440 8352 8492
rect 9680 8440 9732 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10784 8440 10836 8492
rect 7012 8372 7064 8424
rect 11612 8440 11664 8492
rect 12900 8440 12952 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 13912 8372 13964 8424
rect 14188 8372 14240 8424
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 5632 8236 5684 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 8944 8304 8996 8356
rect 10508 8304 10560 8356
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 11152 8304 11204 8356
rect 5908 8236 5960 8245
rect 8208 8236 8260 8288
rect 8760 8236 8812 8288
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 9680 8236 9732 8288
rect 10784 8236 10836 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 13544 8304 13596 8356
rect 12164 8236 12216 8288
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 2412 7828 2464 7880
rect 2504 7828 2556 7880
rect 4160 8032 4212 8084
rect 4344 8032 4396 8084
rect 4988 8032 5040 8084
rect 3884 7896 3936 7948
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 3424 7828 3476 7880
rect 4068 7828 4120 7880
rect 4620 7828 4672 7880
rect 6920 7964 6972 8016
rect 7104 8032 7156 8084
rect 8576 8032 8628 8084
rect 8852 8032 8904 8084
rect 9312 8032 9364 8084
rect 11888 8032 11940 8084
rect 14096 8032 14148 8084
rect 10048 7964 10100 8016
rect 5448 7828 5500 7880
rect 1584 7692 1636 7744
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 4712 7692 4764 7744
rect 6644 7896 6696 7948
rect 9220 7896 9272 7948
rect 9956 7896 10008 7948
rect 13820 7896 13872 7948
rect 7288 7828 7340 7880
rect 7380 7828 7432 7880
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8944 7828 8996 7880
rect 9128 7828 9180 7880
rect 9588 7828 9640 7880
rect 11612 7828 11664 7880
rect 12808 7828 12860 7880
rect 13912 7828 13964 7880
rect 7104 7760 7156 7812
rect 8484 7760 8536 7812
rect 7656 7692 7708 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 8760 7692 8812 7744
rect 9404 7692 9456 7744
rect 12716 7760 12768 7812
rect 13452 7760 13504 7812
rect 13544 7760 13596 7812
rect 11060 7692 11112 7744
rect 12624 7692 12676 7744
rect 12808 7692 12860 7744
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 2136 7488 2188 7540
rect 8392 7488 8444 7540
rect 9588 7488 9640 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 3332 7420 3384 7472
rect 3884 7420 3936 7472
rect 1400 7284 1452 7336
rect 2504 7352 2556 7404
rect 3056 7352 3108 7404
rect 3976 7352 4028 7404
rect 4712 7420 4764 7472
rect 5724 7420 5776 7472
rect 7288 7463 7340 7472
rect 7288 7429 7297 7463
rect 7297 7429 7331 7463
rect 7331 7429 7340 7463
rect 7288 7420 7340 7429
rect 7380 7420 7432 7472
rect 8208 7420 8260 7472
rect 13452 7420 13504 7472
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 3148 7216 3200 7268
rect 3792 7216 3844 7268
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 4988 7216 5040 7268
rect 10232 7352 10284 7404
rect 13912 7488 13964 7540
rect 6000 7216 6052 7268
rect 8300 7284 8352 7336
rect 8392 7284 8444 7336
rect 5264 7148 5316 7200
rect 6644 7148 6696 7200
rect 7104 7148 7156 7200
rect 8300 7148 8352 7200
rect 9956 7148 10008 7200
rect 10968 7148 11020 7200
rect 12808 7284 12860 7336
rect 11704 7216 11756 7268
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 11888 7148 11940 7200
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 3056 6944 3108 6996
rect 5264 6944 5316 6996
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 5632 6944 5684 6996
rect 6184 6944 6236 6996
rect 6552 6944 6604 6996
rect 7012 6944 7064 6996
rect 8944 6944 8996 6996
rect 9496 6944 9548 6996
rect 11612 6944 11664 6996
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2780 6740 2832 6792
rect 3884 6740 3936 6792
rect 4068 6783 4120 6792
rect 4068 6749 4102 6783
rect 4102 6749 4120 6783
rect 4068 6740 4120 6749
rect 3424 6604 3476 6656
rect 4988 6808 5040 6860
rect 7104 6876 7156 6928
rect 5448 6740 5500 6792
rect 8392 6740 8444 6792
rect 5264 6604 5316 6656
rect 7656 6715 7708 6724
rect 7656 6681 7690 6715
rect 7690 6681 7708 6715
rect 7656 6672 7708 6681
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 10416 6808 10468 6860
rect 8760 6604 8812 6613
rect 8944 6604 8996 6656
rect 9220 6672 9272 6724
rect 10232 6672 10284 6724
rect 11612 6808 11664 6860
rect 11888 6808 11940 6860
rect 11704 6672 11756 6724
rect 13268 6740 13320 6792
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 12624 6672 12676 6724
rect 13084 6672 13136 6724
rect 14280 6944 14332 6996
rect 13544 6876 13596 6928
rect 13728 6876 13780 6928
rect 13820 6808 13872 6860
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14004 6740 14056 6792
rect 13820 6604 13872 6656
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2412 6400 2464 6452
rect 3976 6400 4028 6452
rect 5080 6400 5132 6452
rect 5816 6400 5868 6452
rect 5908 6400 5960 6452
rect 7380 6400 7432 6452
rect 7748 6400 7800 6452
rect 8484 6400 8536 6452
rect 2228 6264 2280 6316
rect 2780 6264 2832 6316
rect 3700 6264 3752 6316
rect 4804 6264 4856 6316
rect 7196 6332 7248 6384
rect 3332 6128 3384 6180
rect 3884 6196 3936 6248
rect 3976 6128 4028 6180
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 5448 6196 5500 6248
rect 5632 6128 5684 6180
rect 3884 6060 3936 6112
rect 4068 6060 4120 6112
rect 4344 6060 4396 6112
rect 7380 6264 7432 6316
rect 6092 6196 6144 6248
rect 6920 6196 6972 6248
rect 7012 6196 7064 6248
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 9864 6400 9916 6452
rect 10968 6400 11020 6452
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9128 6264 9180 6316
rect 8944 6196 8996 6248
rect 6184 6128 6236 6180
rect 10784 6264 10836 6316
rect 11704 6400 11756 6452
rect 11244 6332 11296 6384
rect 13544 6400 13596 6452
rect 14372 6443 14424 6452
rect 14372 6409 14381 6443
rect 14381 6409 14415 6443
rect 14415 6409 14424 6443
rect 14372 6400 14424 6409
rect 10140 6196 10192 6248
rect 12808 6332 12860 6384
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 6092 6060 6144 6112
rect 10508 6128 10560 6180
rect 10692 6128 10744 6180
rect 8300 6060 8352 6112
rect 11888 6196 11940 6248
rect 13084 6196 13136 6248
rect 13820 6196 13872 6248
rect 10968 6128 11020 6180
rect 11704 6128 11756 6180
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 11428 6060 11480 6112
rect 12256 6060 12308 6112
rect 14004 6060 14056 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 1768 5856 1820 5908
rect 3056 5856 3108 5908
rect 3700 5856 3752 5908
rect 3792 5856 3844 5908
rect 5264 5856 5316 5908
rect 6000 5856 6052 5908
rect 6736 5856 6788 5908
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 7472 5856 7524 5908
rect 7840 5856 7892 5908
rect 3884 5788 3936 5840
rect 4712 5788 4764 5840
rect 4804 5831 4856 5840
rect 4804 5797 4813 5831
rect 4813 5797 4847 5831
rect 4847 5797 4856 5831
rect 4804 5788 4856 5797
rect 1952 5720 2004 5772
rect 2044 5763 2096 5772
rect 2044 5729 2053 5763
rect 2053 5729 2087 5763
rect 2087 5729 2096 5763
rect 2044 5720 2096 5729
rect 2688 5720 2740 5772
rect 3424 5720 3476 5772
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 5080 5788 5132 5840
rect 6644 5788 6696 5840
rect 1952 5584 2004 5636
rect 2228 5584 2280 5636
rect 2412 5584 2464 5636
rect 5908 5652 5960 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 7012 5652 7064 5704
rect 7380 5788 7432 5840
rect 7196 5652 7248 5704
rect 5632 5584 5684 5636
rect 6092 5584 6144 5636
rect 7748 5652 7800 5704
rect 8760 5788 8812 5840
rect 10140 5788 10192 5840
rect 10048 5720 10100 5772
rect 8392 5652 8444 5704
rect 3424 5516 3476 5568
rect 3884 5516 3936 5568
rect 4988 5516 5040 5568
rect 5264 5516 5316 5568
rect 9864 5584 9916 5636
rect 7656 5516 7708 5568
rect 10416 5516 10468 5568
rect 10968 5856 11020 5908
rect 11060 5856 11112 5908
rect 11428 5856 11480 5908
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 12256 5856 12308 5908
rect 13452 5856 13504 5908
rect 10968 5652 11020 5704
rect 11980 5720 12032 5772
rect 11980 5584 12032 5636
rect 13912 5788 13964 5840
rect 12624 5652 12676 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 12348 5584 12400 5636
rect 12440 5516 12492 5568
rect 14372 5584 14424 5636
rect 14556 5516 14608 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 1308 5312 1360 5364
rect 1952 5312 2004 5364
rect 3056 5312 3108 5364
rect 4252 5312 4304 5364
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 1768 5244 1820 5296
rect 2504 5244 2556 5296
rect 2228 5176 2280 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 4068 5176 4120 5228
rect 4988 5176 5040 5228
rect 5540 5176 5592 5228
rect 5816 5176 5868 5228
rect 6368 5312 6420 5364
rect 6644 5312 6696 5364
rect 6828 5312 6880 5364
rect 9956 5312 10008 5364
rect 8208 5244 8260 5296
rect 10968 5312 11020 5364
rect 12072 5312 12124 5364
rect 14096 5312 14148 5364
rect 14188 5312 14240 5364
rect 6184 5176 6236 5228
rect 6828 5176 6880 5228
rect 6920 5176 6972 5228
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 3332 5108 3384 5160
rect 3608 5108 3660 5160
rect 4160 5108 4212 5160
rect 1768 5040 1820 5092
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5632 5108 5684 5160
rect 5908 5108 5960 5160
rect 3792 4972 3844 5024
rect 8392 5040 8444 5092
rect 9220 5040 9272 5092
rect 12624 5244 12676 5296
rect 12716 5244 12768 5296
rect 13636 5287 13688 5296
rect 13636 5253 13645 5287
rect 13645 5253 13679 5287
rect 13679 5253 13688 5287
rect 13636 5244 13688 5253
rect 10048 5176 10100 5228
rect 11612 5176 11664 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 13360 5176 13412 5228
rect 11244 5108 11296 5160
rect 11060 5040 11112 5092
rect 11888 5108 11940 5160
rect 8300 4972 8352 5024
rect 9956 4972 10008 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 11796 4972 11848 5024
rect 13452 4972 13504 5024
rect 14372 5040 14424 5092
rect 14188 4972 14240 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 1216 4700 1268 4752
rect 2412 4768 2464 4820
rect 3516 4768 3568 4820
rect 3884 4768 3936 4820
rect 4252 4768 4304 4820
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 5908 4768 5960 4820
rect 6092 4768 6144 4820
rect 6828 4768 6880 4820
rect 3148 4700 3200 4752
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 5080 4700 5132 4752
rect 3976 4564 4028 4616
rect 4068 4564 4120 4616
rect 4252 4564 4304 4616
rect 3332 4428 3384 4480
rect 3700 4496 3752 4548
rect 4896 4564 4948 4616
rect 5080 4564 5132 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 9036 4700 9088 4752
rect 9864 4768 9916 4820
rect 10600 4768 10652 4820
rect 10968 4768 11020 4820
rect 11244 4768 11296 4820
rect 12440 4768 12492 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 8392 4632 8444 4684
rect 8576 4632 8628 4684
rect 9864 4632 9916 4684
rect 10232 4632 10284 4684
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 7012 4496 7064 4548
rect 8392 4496 8444 4548
rect 9220 4564 9272 4616
rect 5816 4428 5868 4480
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 7472 4428 7524 4480
rect 9496 4496 9548 4548
rect 10600 4632 10652 4684
rect 10968 4564 11020 4616
rect 12072 4632 12124 4684
rect 12808 4675 12860 4684
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 11980 4496 12032 4548
rect 13728 4768 13780 4820
rect 13636 4564 13688 4616
rect 13544 4539 13596 4548
rect 13544 4505 13553 4539
rect 13553 4505 13587 4539
rect 13587 4505 13596 4539
rect 13544 4496 13596 4505
rect 13452 4428 13504 4480
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 1768 4267 1820 4276
rect 1768 4233 1777 4267
rect 1777 4233 1811 4267
rect 1811 4233 1820 4267
rect 1768 4224 1820 4233
rect 2228 4224 2280 4276
rect 1584 4088 1636 4140
rect 2504 4156 2556 4208
rect 3700 4267 3752 4276
rect 3700 4233 3709 4267
rect 3709 4233 3743 4267
rect 3743 4233 3752 4267
rect 3700 4224 3752 4233
rect 4804 4224 4856 4276
rect 5540 4224 5592 4276
rect 6092 4224 6144 4276
rect 6368 4224 6420 4276
rect 4344 4156 4396 4208
rect 1032 4020 1084 4072
rect 2964 4088 3016 4140
rect 3516 4088 3568 4140
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 2412 4063 2464 4072
rect 2412 4029 2421 4063
rect 2421 4029 2455 4063
rect 2455 4029 2464 4063
rect 2412 4020 2464 4029
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 3332 4020 3384 4072
rect 4804 4020 4856 4072
rect 6828 4156 6880 4208
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 8300 4224 8352 4276
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 8760 4224 8812 4276
rect 9036 4224 9088 4276
rect 10140 4224 10192 4276
rect 13544 4224 13596 4276
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 7012 4088 7064 4140
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 2504 3884 2556 3936
rect 2872 3884 2924 3936
rect 4620 3952 4672 4004
rect 5724 3952 5776 4004
rect 6552 4020 6604 4072
rect 7104 4020 7156 4072
rect 7196 4020 7248 4072
rect 4804 3884 4856 3936
rect 6276 3884 6328 3936
rect 7104 3884 7156 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7288 3884 7340 3936
rect 7472 3884 7524 3936
rect 7748 4020 7800 4072
rect 7656 3952 7708 4004
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 9864 4156 9916 4208
rect 10600 4156 10652 4208
rect 9404 4088 9456 4140
rect 11428 4156 11480 4208
rect 11244 4088 11296 4140
rect 13084 4088 13136 4140
rect 8576 3952 8628 4004
rect 9036 3884 9088 3936
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 11704 4020 11756 4072
rect 11980 4020 12032 4072
rect 12072 4020 12124 4072
rect 12348 4020 12400 4072
rect 14004 4156 14056 4208
rect 13360 4088 13412 4140
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 11336 3884 11388 3936
rect 11704 3884 11756 3936
rect 12624 3884 12676 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 1124 3680 1176 3732
rect 1860 3680 1912 3732
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2780 3680 2832 3732
rect 3148 3680 3200 3732
rect 3700 3680 3752 3732
rect 4160 3680 4212 3732
rect 4252 3680 4304 3732
rect 6644 3680 6696 3732
rect 7104 3680 7156 3732
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 7840 3680 7892 3732
rect 1584 3612 1636 3664
rect 3792 3612 3844 3664
rect 7472 3612 7524 3664
rect 2780 3476 2832 3528
rect 4252 3544 4304 3596
rect 4712 3544 4764 3596
rect 10416 3612 10468 3664
rect 10600 3612 10652 3664
rect 10692 3655 10744 3664
rect 10692 3621 10701 3655
rect 10701 3621 10735 3655
rect 10735 3621 10744 3655
rect 10692 3612 10744 3621
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11612 3680 11664 3732
rect 12072 3680 12124 3732
rect 14096 3680 14148 3732
rect 8208 3544 8260 3596
rect 8300 3544 8352 3596
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 11888 3587 11940 3596
rect 756 3340 808 3392
rect 3700 3408 3752 3460
rect 4620 3408 4672 3460
rect 4988 3476 5040 3528
rect 9404 3476 9456 3528
rect 10692 3476 10744 3528
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 11612 3476 11664 3528
rect 5816 3408 5868 3460
rect 7012 3408 7064 3460
rect 7104 3408 7156 3460
rect 7840 3340 7892 3392
rect 8576 3408 8628 3460
rect 11888 3408 11940 3460
rect 11980 3408 12032 3460
rect 14372 3544 14424 3596
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 13728 3476 13780 3528
rect 14556 3408 14608 3460
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 2320 3136 2372 3188
rect 3332 3136 3384 3188
rect 4068 3136 4120 3188
rect 4160 3136 4212 3188
rect 5080 3136 5132 3188
rect 6552 3136 6604 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7196 3136 7248 3188
rect 3884 3068 3936 3120
rect 1308 3000 1360 3052
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 480 2932 532 2984
rect 572 2932 624 2984
rect 1492 2907 1544 2916
rect 1492 2873 1501 2907
rect 1501 2873 1535 2907
rect 1535 2873 1544 2907
rect 1492 2864 1544 2873
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 3240 3000 3292 3052
rect 3516 3000 3568 3052
rect 4068 3000 4120 3052
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 6644 3000 6696 3052
rect 6736 3000 6788 3052
rect 2964 2864 3016 2916
rect 5540 2975 5592 2984
rect 5540 2941 5549 2975
rect 5549 2941 5583 2975
rect 5583 2941 5592 2975
rect 5540 2932 5592 2941
rect 6920 3068 6972 3120
rect 7656 3068 7708 3120
rect 8208 3068 8260 3120
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 9036 3136 9088 3188
rect 9588 3136 9640 3188
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 11704 3136 11756 3188
rect 11888 3136 11940 3188
rect 12256 3136 12308 3188
rect 9220 3068 9272 3120
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 8300 3000 8352 3052
rect 13636 3136 13688 3188
rect 3976 2864 4028 2916
rect 4344 2796 4396 2848
rect 5540 2796 5592 2848
rect 7012 2864 7064 2916
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 7380 2932 7432 2984
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 9588 2932 9640 2984
rect 9220 2864 9272 2916
rect 10692 3000 10744 3052
rect 12532 3068 12584 3120
rect 13360 3068 13412 3120
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 7932 2796 7984 2848
rect 9404 2796 9456 2848
rect 10876 2932 10928 2984
rect 12164 2932 12216 2984
rect 12716 2932 12768 2984
rect 14464 3000 14516 3052
rect 14372 2932 14424 2984
rect 11612 2864 11664 2916
rect 13820 2864 13872 2916
rect 10140 2796 10192 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 388 2592 440 2644
rect 2504 2592 2556 2644
rect 3056 2592 3108 2644
rect 664 2524 716 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 5080 2592 5132 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 7840 2592 7892 2644
rect 9680 2592 9732 2644
rect 10508 2592 10560 2644
rect 12808 2592 12860 2644
rect 4804 2524 4856 2576
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2228 2388 2280 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 3240 2388 3292 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 3700 2320 3752 2372
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5448 2456 5500 2508
rect 5540 2456 5592 2508
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 8116 2456 8168 2508
rect 5264 2388 5316 2440
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 5632 2388 5684 2440
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 4528 2252 4580 2304
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 5264 2252 5316 2304
rect 6644 2252 6696 2304
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 7104 2363 7156 2372
rect 7104 2329 7113 2363
rect 7113 2329 7147 2363
rect 7147 2329 7156 2363
rect 7104 2320 7156 2329
rect 7196 2320 7248 2372
rect 8576 2524 8628 2576
rect 9772 2456 9824 2508
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 8576 2320 8628 2372
rect 9404 2320 9456 2372
rect 8668 2252 8720 2304
rect 11980 2524 12032 2576
rect 10324 2456 10376 2508
rect 10784 2456 10836 2508
rect 13360 2524 13412 2576
rect 14280 2592 14332 2644
rect 12808 2456 12860 2508
rect 13268 2499 13320 2508
rect 13268 2465 13277 2499
rect 13277 2465 13311 2499
rect 13311 2465 13320 2499
rect 13268 2456 13320 2465
rect 10416 2388 10468 2440
rect 11152 2388 11204 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 11704 2363 11756 2372
rect 11704 2329 11713 2363
rect 11713 2329 11747 2363
rect 11747 2329 11756 2363
rect 11704 2320 11756 2329
rect 11888 2320 11940 2372
rect 12440 2363 12492 2372
rect 12440 2329 12449 2363
rect 12449 2329 12483 2363
rect 12483 2329 12492 2363
rect 12440 2320 12492 2329
rect 12532 2363 12584 2372
rect 12532 2329 12541 2363
rect 12541 2329 12575 2363
rect 12575 2329 12584 2363
rect 12532 2320 12584 2329
rect 10968 2252 11020 2304
rect 12164 2252 12216 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 1676 2048 1728 2100
rect 2412 2048 2464 2100
rect 3792 2048 3844 2100
rect 6736 2048 6788 2100
rect 13084 2048 13136 2100
rect 4896 1980 4948 2032
rect 8300 1980 8352 2032
rect 8484 1980 8536 2032
rect 8760 1980 8812 2032
rect 9956 1980 10008 2032
rect 12164 1980 12216 2032
rect 4712 1912 4764 1964
rect 11152 1912 11204 1964
rect 4804 1844 4856 1896
rect 12716 1844 12768 1896
rect 2964 1776 3016 1828
rect 7196 1776 7248 1828
rect 3976 1708 4028 1760
rect 9772 1776 9824 1828
rect 8208 1708 8260 1760
rect 11244 1708 11296 1760
rect 8944 1640 8996 1692
rect 4988 1300 5040 1352
rect 9956 1300 10008 1352
rect 10232 1232 10284 1284
rect 12348 1232 12400 1284
<< metal2 >>
rect 2778 18592 2834 18601
rect 2778 18527 2834 18536
rect 13726 18592 13782 18601
rect 13726 18527 13782 18536
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 952 16794 980 17711
rect 2792 17270 2820 18527
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 13740 17338 13768 18527
rect 14646 17776 14702 17785
rect 14568 17734 14646 17762
rect 14568 17338 14596 17734
rect 14646 17711 14702 17720
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 1032 16992 1084 16998
rect 1030 16960 1032 16969
rect 1084 16960 1086 16969
rect 1030 16895 1086 16904
rect 2424 16794 2452 17138
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 940 16788 992 16794
rect 940 16730 992 16736
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 940 16244 992 16250
rect 940 16186 992 16192
rect 952 16153 980 16186
rect 938 16144 994 16153
rect 938 16079 994 16088
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 1136 15337 1164 15642
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 1584 15360 1636 15366
rect 1122 15328 1178 15337
rect 1584 15302 1636 15308
rect 1122 15263 1178 15272
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 14618 1440 14758
rect 1596 14657 1624 15302
rect 2884 15026 2912 15370
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 1582 14648 1638 14657
rect 1400 14612 1452 14618
rect 1582 14583 1638 14592
rect 1400 14554 1452 14560
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1216 14068 1268 14074
rect 1216 14010 1268 14016
rect 480 13932 532 13938
rect 480 13874 532 13880
rect 388 12912 440 12918
rect 388 12854 440 12860
rect 400 2650 428 12854
rect 492 2990 520 13874
rect 756 13796 808 13802
rect 756 13738 808 13744
rect 572 13388 624 13394
rect 572 13330 624 13336
rect 584 3369 612 13330
rect 664 13252 716 13258
rect 664 13194 716 13200
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 388 2644 440 2650
rect 388 2586 440 2592
rect 584 800 612 2926
rect 676 2582 704 13194
rect 768 3398 796 13738
rect 1124 13456 1176 13462
rect 1124 13398 1176 13404
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 952 12889 980 13126
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 848 12640 900 12646
rect 848 12582 900 12588
rect 756 3392 808 3398
rect 756 3334 808 3340
rect 664 2576 716 2582
rect 664 2518 716 2524
rect 570 0 626 800
rect 860 762 888 12582
rect 1030 12336 1086 12345
rect 1030 12271 1086 12280
rect 940 12096 992 12102
rect 938 12064 940 12073
rect 992 12064 994 12073
rect 938 11999 994 12008
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10441 980 10610
rect 938 10432 994 10441
rect 938 10367 994 10376
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 952 8974 980 9551
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 952 4729 980 8774
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1044 4078 1072 12271
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 1136 3738 1164 13398
rect 1228 12434 1256 14010
rect 1504 14006 1532 14311
rect 1688 14006 1716 14962
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1872 14278 1900 14350
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1492 14000 1544 14006
rect 1492 13942 1544 13948
rect 1676 14000 1728 14006
rect 1676 13942 1728 13948
rect 1584 13728 1636 13734
rect 1582 13696 1584 13705
rect 1636 13696 1638 13705
rect 1582 13631 1638 13640
rect 1584 12640 1636 12646
rect 1582 12608 1584 12617
rect 1636 12608 1638 12617
rect 1582 12543 1638 12552
rect 1228 12406 1348 12434
rect 1216 11620 1268 11626
rect 1216 11562 1268 11568
rect 1228 4758 1256 11562
rect 1320 5370 1348 12406
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1504 11898 1532 12106
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1688 11762 1716 13942
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1688 11558 1716 11698
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1412 10554 1440 11494
rect 1492 11348 1544 11354
rect 1780 11336 1808 12786
rect 1544 11308 1808 11336
rect 1492 11290 1544 11296
rect 1676 11144 1728 11150
rect 1674 11112 1676 11121
rect 1728 11112 1730 11121
rect 1674 11047 1730 11056
rect 1872 10713 1900 14214
rect 1964 12434 1992 14758
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2410 14512 2466 14521
rect 2410 14447 2412 14456
rect 2464 14447 2466 14456
rect 2412 14418 2464 14424
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2976 14226 3004 14350
rect 3252 14249 3280 14758
rect 3344 14278 3372 14758
rect 3332 14272 3384 14278
rect 3238 14240 3294 14249
rect 2056 12850 2084 14214
rect 2976 14198 3188 14226
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2332 13841 2360 13874
rect 2318 13832 2374 13841
rect 2318 13767 2374 13776
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 12986 2176 13262
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1964 12406 2268 12434
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 11665 2084 11698
rect 2042 11656 2098 11665
rect 2042 11591 2098 11600
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1858 10704 1914 10713
rect 1858 10639 1914 10648
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1676 10600 1728 10606
rect 1412 10526 1532 10554
rect 1676 10542 1728 10548
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9722 1440 10406
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 7886 1440 8774
rect 1504 7993 1532 10526
rect 1688 9722 1716 10542
rect 1964 9722 1992 10610
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 8430 1716 9454
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 8498 1808 9318
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1858 8392 1914 8401
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1490 7848 1546 7857
rect 1490 7783 1492 7792
rect 1544 7783 1546 7792
rect 1492 7754 1544 7760
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1490 7304 1546 7313
rect 1412 6798 1440 7278
rect 1490 7239 1546 7248
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1216 4752 1268 4758
rect 1216 4694 1268 4700
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1320 3058 1348 5199
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1412 2514 1440 6287
rect 1504 4026 1532 7239
rect 1596 4146 1624 7686
rect 1688 5794 1716 8366
rect 1768 8356 1820 8362
rect 1858 8327 1914 8336
rect 1768 8298 1820 8304
rect 1780 7562 1808 8298
rect 1872 7886 1900 8327
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1780 7534 1900 7562
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 5914 1808 7346
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1688 5766 1808 5794
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1504 3998 1624 4026
rect 1596 3670 1624 3998
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1688 3058 1716 5471
rect 1780 5302 1808 5766
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 1780 4282 1808 5034
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1872 3738 1900 7534
rect 2056 6984 2084 11086
rect 2148 10452 2176 11494
rect 2240 10554 2268 12406
rect 2332 10849 2360 13126
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 11694 2452 12582
rect 2516 12442 2544 13874
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2976 12850 3004 13194
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2962 12744 3018 12753
rect 2962 12679 2964 12688
rect 3016 12679 3018 12688
rect 2964 12650 3016 12656
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2516 11558 2544 12106
rect 2884 11898 2912 12106
rect 3068 12073 3096 14010
rect 3160 13274 3188 14198
rect 3332 14214 3384 14220
rect 3238 14175 3294 14184
rect 3436 14074 3464 15438
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3528 14414 3556 14554
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3528 13920 3556 14214
rect 3436 13892 3556 13920
rect 3436 13802 3464 13892
rect 3620 13818 3648 14826
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3712 14074 3740 14418
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3804 14006 3832 14282
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3792 13864 3844 13870
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3516 13796 3568 13802
rect 3620 13790 3740 13818
rect 4080 13841 4108 13874
rect 3792 13806 3844 13812
rect 4066 13832 4122 13841
rect 3516 13738 3568 13744
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3252 13394 3280 13670
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3344 13326 3372 13670
rect 3332 13320 3384 13326
rect 3238 13288 3294 13297
rect 3160 13246 3238 13274
rect 3332 13262 3384 13268
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3238 13223 3294 13232
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 13025 3372 13126
rect 3330 13016 3386 13025
rect 3330 12951 3386 12960
rect 3240 12640 3292 12646
rect 3238 12608 3240 12617
rect 3436 12628 3464 13262
rect 3292 12608 3294 12617
rect 3238 12543 3294 12552
rect 3344 12600 3464 12628
rect 3240 12096 3292 12102
rect 3054 12064 3110 12073
rect 3240 12038 3292 12044
rect 3054 11999 3110 12008
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11336 2544 11494
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 3160 11354 3188 11698
rect 3148 11348 3200 11354
rect 2516 11308 2820 11336
rect 2792 11150 2820 11308
rect 3148 11290 3200 11296
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3054 11112 3110 11121
rect 3054 11047 3110 11056
rect 3068 11014 3096 11047
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2318 10840 2374 10849
rect 2318 10775 2374 10784
rect 3160 10674 3188 10950
rect 3252 10674 3280 12038
rect 3344 10810 3372 12600
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 12102 3464 12378
rect 3528 12306 3556 13738
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3620 12186 3648 13126
rect 3528 12158 3648 12186
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11354 3464 11766
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 2318 10568 2374 10577
rect 2240 10526 2318 10554
rect 2318 10503 2374 10512
rect 2148 10424 2268 10452
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 2148 8634 2176 9930
rect 2240 9081 2268 10424
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9586 3096 9998
rect 3160 9722 3188 10610
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2226 9072 2282 9081
rect 2226 9007 2282 9016
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 7546 2176 8366
rect 2240 8090 2268 8910
rect 2332 8838 2360 9415
rect 2424 9178 2452 9522
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2318 7984 2374 7993
rect 2240 7942 2318 7970
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1964 6956 2084 6984
rect 1964 5778 1992 6956
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 2056 5778 2084 6831
rect 2240 6474 2268 7942
rect 2318 7919 2374 7928
rect 2424 7886 2452 8774
rect 2504 8424 2556 8430
rect 2608 8401 2636 8910
rect 2700 8498 2728 9114
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 3068 8430 3096 9522
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 9178 3188 9454
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3056 8424 3108 8430
rect 2504 8366 2556 8372
rect 2594 8392 2650 8401
rect 2516 7886 2544 8366
rect 3056 8366 3108 8372
rect 2594 8327 2650 8336
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 3068 7410 3096 8366
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2240 6446 2360 6474
rect 2424 6458 2452 7142
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2240 5642 2268 6258
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 1964 5370 1992 5578
rect 2332 5386 2360 6446
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2056 5358 2360 5386
rect 1950 4584 2006 4593
rect 1950 4519 2006 4528
rect 1964 3942 1992 4519
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1490 2952 1546 2961
rect 1490 2887 1492 2896
rect 1544 2887 1546 2896
rect 1492 2858 1544 2864
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 2106 1716 2382
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1228 870 1348 898
rect 1228 762 1256 870
rect 1320 800 1348 870
rect 2056 800 2084 5358
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2240 4282 2268 5170
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2240 2446 2268 4111
rect 2332 3194 2360 5170
rect 2424 4826 2452 5578
rect 2516 5302 2544 7346
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 3068 7002 3096 7346
rect 3160 7274 3188 8842
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6322 2820 6734
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 3068 5914 3096 6938
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2700 5148 2728 5714
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2516 5120 2728 5148
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2516 4214 2544 5120
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2412 4072 2464 4078
rect 2410 4040 2412 4049
rect 2464 4040 2466 4049
rect 2410 3975 2466 3984
rect 2884 3942 2912 4558
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2976 4049 3004 4082
rect 2962 4040 3018 4049
rect 2962 3975 3018 3984
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2516 3738 2544 3878
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2792 3534 2820 3674
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2700 2922 3004 2938
rect 2700 2916 3016 2922
rect 2700 2910 2964 2916
rect 2412 2848 2464 2854
rect 2700 2836 2728 2910
rect 2964 2858 3016 2864
rect 2412 2790 2464 2796
rect 2516 2808 2728 2836
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2424 2106 2452 2790
rect 2516 2650 2544 2808
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 3068 2650 3096 5306
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3160 3738 3188 4694
rect 3252 4162 3280 10406
rect 3344 7478 3372 10542
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 10198 3464 10406
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3424 9920 3476 9926
rect 3422 9888 3424 9897
rect 3476 9888 3478 9897
rect 3422 9823 3478 9832
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9353 3464 9522
rect 3422 9344 3478 9353
rect 3422 9279 3478 9288
rect 3436 9110 3464 9279
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3344 6186 3372 7414
rect 3436 6662 3464 7822
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3436 5778 3464 6598
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3424 5568 3476 5574
rect 3528 5556 3556 12158
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11286 3648 12038
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 9926 3648 10950
rect 3712 10062 3740 13790
rect 3804 12209 3832 13806
rect 4066 13767 4122 13776
rect 4172 12782 4200 14894
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 13841 4752 13874
rect 4710 13832 4766 13841
rect 4710 13767 4766 13776
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3896 12424 3924 12543
rect 4080 12442 4108 12718
rect 4068 12436 4120 12442
rect 3896 12396 4016 12424
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11898 3832 12038
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3896 11778 3924 12242
rect 3804 11750 3924 11778
rect 3804 10849 3832 11750
rect 3988 11642 4016 12396
rect 4068 12378 4120 12384
rect 4172 12374 4200 12718
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3896 11614 4016 11642
rect 3790 10840 3846 10849
rect 3790 10775 3846 10784
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3804 10266 3832 10610
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 8566 3648 9862
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3712 8378 3740 9658
rect 3804 8498 3832 10202
rect 3896 10062 3924 11614
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11098 4016 11494
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4080 11257 4108 11290
rect 4066 11248 4122 11257
rect 4066 11183 4122 11192
rect 4068 11144 4120 11150
rect 3988 11092 4068 11098
rect 3988 11086 4120 11092
rect 3988 11070 4108 11086
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10470 4016 10950
rect 4080 10810 4108 11070
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10266 4016 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3896 9722 3924 9998
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3476 5528 3556 5556
rect 3620 8350 3740 8378
rect 3424 5510 3476 5516
rect 3620 5166 3648 8350
rect 3804 7274 3832 8434
rect 3988 8362 4016 9114
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3896 7954 3924 8298
rect 4080 8072 4108 10639
rect 4172 8634 4200 12106
rect 4264 11898 4292 12854
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4356 12306 4384 12718
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4540 12170 4568 12854
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4632 12434 4660 12786
rect 4632 12406 4752 12434
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4724 12102 4752 12406
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4724 11762 4752 12038
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4250 11656 4306 11665
rect 4724 11626 4752 11698
rect 4250 11591 4306 11600
rect 4712 11620 4764 11626
rect 4264 11082 4292 11591
rect 4712 11562 4764 11568
rect 4816 11200 4844 13942
rect 4724 11172 4844 11200
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4264 9722 4292 9998
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4264 9178 4292 9658
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4724 9081 4752 11172
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4710 9072 4766 9081
rect 4710 9007 4766 9016
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4172 8090 4200 8570
rect 3988 8044 4108 8072
rect 4160 8084 4212 8090
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3884 7744 3936 7750
rect 3988 7721 4016 8044
rect 4160 8026 4212 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3884 7686 3936 7692
rect 3974 7712 4030 7721
rect 3896 7478 3924 7686
rect 3974 7647 4030 7656
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3882 7032 3938 7041
rect 3804 6990 3882 7018
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3712 5914 3740 6258
rect 3804 5914 3832 6990
rect 3882 6967 3938 6976
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6254 3924 6734
rect 3988 6458 4016 7346
rect 4080 6798 4108 7822
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3988 6186 4200 6202
rect 3976 6180 4200 6186
rect 4028 6174 4200 6180
rect 3976 6122 4028 6128
rect 3884 6112 3936 6118
rect 4068 6112 4120 6118
rect 3884 6054 3936 6060
rect 3974 6080 4030 6089
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3896 5846 3924 6054
rect 4068 6054 4120 6060
rect 3974 6015 4030 6024
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3332 5160 3384 5166
rect 3608 5160 3660 5166
rect 3514 5128 3570 5137
rect 3332 5102 3384 5108
rect 3344 4486 3372 5102
rect 3436 5086 3514 5114
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3252 4134 3372 4162
rect 3344 4078 3372 4134
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3160 2774 3188 3674
rect 3252 3505 3280 4014
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 3238 3360 3294 3369
rect 3238 3295 3294 3304
rect 3252 3058 3280 3295
rect 3344 3194 3372 3839
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3436 2904 3464 5086
rect 3608 5102 3660 5108
rect 3514 5063 3570 5072
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3528 4146 3556 4762
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4282 3740 4490
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3528 3058 3556 4082
rect 3712 3738 3740 4218
rect 3804 4146 3832 4966
rect 3896 4826 3924 5510
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3988 4706 4016 6015
rect 4080 5234 4108 6054
rect 4172 5250 4200 6174
rect 4264 5710 4292 8774
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4724 8537 4752 8910
rect 4710 8528 4766 8537
rect 4620 8492 4672 8498
rect 4710 8463 4766 8472
rect 4620 8434 4672 8440
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 8090 4384 8230
rect 4434 8120 4490 8129
rect 4344 8084 4396 8090
rect 4434 8055 4490 8064
rect 4344 8026 4396 8032
rect 4448 7954 4476 8055
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4632 7886 4660 8434
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 4724 7478 4752 7686
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 4816 6440 4844 11018
rect 4908 10305 4936 14962
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 5000 13025 5028 13126
rect 4986 13016 5042 13025
rect 4986 12951 5042 12960
rect 5092 12434 5120 14010
rect 5172 13184 5224 13190
rect 5276 13161 5304 14214
rect 5172 13126 5224 13132
rect 5262 13152 5318 13161
rect 5184 12889 5212 13126
rect 5262 13087 5318 13096
rect 5170 12880 5226 12889
rect 5170 12815 5226 12824
rect 5264 12776 5316 12782
rect 5538 12744 5594 12753
rect 5264 12718 5316 12724
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5000 12406 5120 12434
rect 4894 10296 4950 10305
rect 4894 10231 4950 10240
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4724 6412 4844 6440
rect 4618 6352 4674 6361
rect 4618 6287 4674 6296
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4356 5556 4384 6054
rect 4264 5528 4384 5556
rect 4632 5556 4660 6287
rect 4724 5846 4752 6412
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4816 5846 4844 6258
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4632 5528 4752 5556
rect 4264 5370 4292 5528
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4068 5228 4120 5234
rect 4172 5222 4292 5250
rect 4068 5170 4120 5176
rect 3896 4678 4016 4706
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3790 3768 3846 3777
rect 3700 3732 3752 3738
rect 3790 3703 3846 3712
rect 3700 3674 3752 3680
rect 3804 3670 3832 3703
rect 3792 3664 3844 3670
rect 3896 3641 3924 4678
rect 4080 4622 4108 5170
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3792 3606 3844 3612
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 3882 3496 3938 3505
rect 3700 3460 3752 3466
rect 3882 3431 3938 3440
rect 3700 3402 3752 3408
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3436 2876 3556 2904
rect 3160 2746 3280 2774
rect 3146 2680 3202 2689
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 3056 2644 3108 2650
rect 3146 2615 3202 2624
rect 3056 2586 3108 2592
rect 2594 2544 2650 2553
rect 2594 2479 2650 2488
rect 2608 2446 2636 2479
rect 3160 2446 3188 2615
rect 3252 2446 3280 2746
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3344 2310 3372 2343
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 2976 1834 3004 2246
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 2700 870 2820 898
rect 860 734 1256 762
rect 1306 0 1362 800
rect 2042 0 2098 800
rect 2700 785 2728 870
rect 2792 800 2820 870
rect 3528 800 3556 2876
rect 3712 2378 3740 3402
rect 3896 3126 3924 3431
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3988 2922 4016 4558
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4080 3194 4108 4111
rect 4172 3738 4200 5102
rect 4264 4826 4292 5222
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 3738 4292 4558
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4172 3194 4200 3674
rect 4252 3596 4304 3602
rect 4356 3584 4384 4150
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4304 3556 4384 3584
rect 4252 3538 4304 3544
rect 4632 3466 4660 3946
rect 4724 3602 4752 5528
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4282 4844 4762
rect 4908 4622 4936 10134
rect 5000 8634 5028 12406
rect 5184 12345 5212 12582
rect 5170 12336 5226 12345
rect 5170 12271 5226 12280
rect 5276 12220 5304 12718
rect 5092 12192 5304 12220
rect 5460 12702 5538 12730
rect 5092 9382 5120 12192
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 11898 5396 12106
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5262 11792 5318 11801
rect 5262 11727 5318 11736
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 10810 5212 11630
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5184 9722 5212 10746
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 7274 5028 8026
rect 5092 7449 5120 8910
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5078 7440 5134 7449
rect 5078 7375 5134 7384
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 5658 5028 6802
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5092 5846 5120 6394
rect 5184 6089 5212 8842
rect 5276 8276 5304 11727
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 8566 5396 9862
rect 5460 9674 5488 12702
rect 5538 12679 5594 12688
rect 5644 12434 5672 17070
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5736 12617 5764 12786
rect 5816 12776 5868 12782
rect 5814 12744 5816 12753
rect 5868 12744 5870 12753
rect 5814 12679 5870 12688
rect 5722 12608 5778 12617
rect 5722 12543 5778 12552
rect 5644 12406 5856 12434
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11150 5580 12174
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10470 5580 10950
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 9994 5580 10406
rect 5644 10305 5672 12038
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11286 5764 11494
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5460 9646 5580 9674
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5276 8248 5396 8276
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 7002 5304 7142
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5170 6080 5226 6089
rect 5170 6015 5226 6024
rect 5276 5914 5304 6598
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5000 5630 5120 5658
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 5234 5028 5510
rect 5092 5370 5120 5630
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5078 5264 5134 5273
rect 4988 5228 5040 5234
rect 5134 5222 5212 5250
rect 5078 5199 5134 5208
rect 4988 5170 5040 5176
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4894 4448 4950 4457
rect 4894 4383 4950 4392
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4804 4072 4856 4078
rect 4802 4040 4804 4049
rect 4856 4040 4858 4049
rect 4802 3975 4858 3984
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4816 3058 4844 3878
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4080 2553 4108 2994
rect 4908 2938 4936 4383
rect 5000 3534 5028 5170
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5092 4622 5120 4694
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5092 3194 5120 4558
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4986 3088 5042 3097
rect 4986 3023 4988 3032
rect 5040 3023 5042 3032
rect 4988 2994 5040 3000
rect 4632 2910 4936 2938
rect 4344 2848 4396 2854
rect 4250 2816 4306 2825
rect 4344 2790 4396 2796
rect 4250 2751 4306 2760
rect 4066 2544 4122 2553
rect 4066 2479 4122 2488
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3804 2106 3832 2382
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3988 1766 4016 2246
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 4264 800 4292 2751
rect 4356 2446 4384 2790
rect 4632 2774 4660 2910
rect 5184 2774 5212 5222
rect 5276 3913 5304 5510
rect 5368 5166 5396 8248
rect 5460 7993 5488 8774
rect 5446 7984 5502 7993
rect 5446 7919 5502 7928
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7002 5488 7822
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6254 5488 6734
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5552 5522 5580 9646
rect 5630 9344 5686 9353
rect 5630 9279 5686 9288
rect 5644 8974 5672 9279
rect 5736 9178 5764 9998
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 7002 5672 8230
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5736 6202 5764 7414
rect 5828 6882 5856 12406
rect 5920 10112 5948 15302
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12238 6040 13194
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6012 10810 6040 11698
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6564 11286 6592 11630
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6012 10266 6040 10474
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6000 10124 6052 10130
rect 5920 10084 6000 10112
rect 6000 10066 6052 10072
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9674 6040 9862
rect 5920 9646 6040 9674
rect 5920 9518 5948 9646
rect 6000 9580 6052 9586
rect 6104 9568 6132 10066
rect 6196 9722 6224 10202
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6380 9586 6408 10134
rect 6472 9722 6500 10542
rect 6564 10266 6592 10678
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6550 10160 6606 10169
rect 6550 10095 6606 10104
rect 6564 9722 6592 10095
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6052 9540 6132 9568
rect 6368 9580 6420 9586
rect 6000 9522 6052 9528
rect 6368 9522 6420 9528
rect 5908 9512 5960 9518
rect 6656 9500 6684 12582
rect 6748 12306 6776 12718
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11830 6868 12174
rect 6828 11824 6880 11830
rect 6932 11801 6960 13806
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 6828 11766 6880 11772
rect 6918 11792 6974 11801
rect 6918 11727 6974 11736
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6840 11082 6868 11562
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 9926 6776 10406
rect 6932 10130 6960 11630
rect 7116 11257 7144 12854
rect 7208 12306 7236 15030
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12442 7328 12786
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7668 11830 7696 13806
rect 8128 13530 8156 13806
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11286 7328 11494
rect 7484 11354 7512 11698
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7288 11280 7340 11286
rect 7102 11248 7158 11257
rect 7288 11222 7340 11228
rect 7102 11183 7158 11192
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10810 7144 11018
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9654 6776 9862
rect 7116 9738 7144 10474
rect 7024 9710 7144 9738
rect 7024 9674 7052 9710
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 9646 7052 9674
rect 7104 9648 7156 9654
rect 6736 9512 6788 9518
rect 5908 9454 5960 9460
rect 6472 9472 6736 9500
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8294 5948 9318
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 8129 5948 8230
rect 5906 8120 5962 8129
rect 5906 8055 5962 8064
rect 6012 7410 6040 9046
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 8634 6316 8910
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8276 6408 8774
rect 6472 8566 6500 9472
rect 6736 9454 6788 9460
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6564 8906 6592 9318
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6564 8498 6592 8842
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 8424 6512 8430
rect 6512 8372 6592 8378
rect 6460 8366 6592 8372
rect 6472 8350 6592 8366
rect 6380 8248 6500 8276
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5828 6854 5948 6882
rect 5920 6458 5948 6854
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5644 6186 5764 6202
rect 5632 6180 5764 6186
rect 5684 6174 5764 6180
rect 5828 6202 5856 6394
rect 5908 6316 5960 6322
rect 6012 6304 6040 7210
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 5960 6276 6040 6304
rect 5908 6258 5960 6264
rect 6092 6248 6144 6254
rect 5828 6196 6092 6202
rect 5828 6190 6144 6196
rect 5828 6174 6132 6190
rect 6196 6186 6224 6938
rect 6184 6180 6236 6186
rect 5632 6122 5684 6128
rect 6184 6122 6236 6128
rect 6092 6112 6144 6118
rect 5920 6072 6092 6100
rect 5920 5710 5948 6072
rect 6092 6054 6144 6060
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5908 5704 5960 5710
rect 5814 5672 5870 5681
rect 5632 5636 5684 5642
rect 5908 5646 5960 5652
rect 5814 5607 5870 5616
rect 5632 5578 5684 5584
rect 5460 5494 5580 5522
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5354 4720 5410 4729
rect 5354 4655 5410 4664
rect 5368 4622 5396 4655
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 4540 2746 4660 2774
rect 5092 2746 5212 2774
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4540 2310 4568 2746
rect 4618 2680 4674 2689
rect 5092 2650 5120 2746
rect 4618 2615 4674 2624
rect 5080 2644 5132 2650
rect 4632 2446 4660 2615
rect 5080 2586 5132 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 4724 1970 4752 2246
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4816 1902 4844 2518
rect 5460 2514 5488 5494
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5552 4826 5580 5170
rect 5644 5166 5672 5578
rect 5828 5234 5856 5607
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5552 4282 5580 4762
rect 6012 4622 6040 5850
rect 6366 5808 6422 5817
rect 6366 5743 6422 5752
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5137 6132 5578
rect 6182 5400 6238 5409
rect 6380 5370 6408 5743
rect 6182 5335 6238 5344
rect 6368 5364 6420 5370
rect 6196 5234 6224 5335
rect 6368 5306 6420 5312
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6090 5128 6146 5137
rect 6090 5063 6146 5072
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6000 4616 6052 4622
rect 5920 4576 6000 4604
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5722 4312 5778 4321
rect 5540 4276 5592 4282
rect 5722 4247 5778 4256
rect 5540 4218 5592 4224
rect 5736 4010 5764 4247
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5722 3768 5778 3777
rect 5722 3703 5778 3712
rect 5630 3632 5686 3641
rect 5630 3567 5686 3576
rect 5644 3210 5672 3567
rect 5736 3369 5764 3703
rect 5828 3466 5856 4422
rect 5920 4146 5948 4576
rect 6000 4558 6052 4564
rect 6104 4282 6132 4762
rect 6366 4312 6422 4321
rect 6092 4276 6144 4282
rect 6366 4247 6368 4256
rect 6092 4218 6144 4224
rect 6420 4247 6422 4256
rect 6368 4218 6420 4224
rect 6472 4162 6500 8248
rect 6564 7188 6592 8350
rect 6656 7954 6684 8978
rect 6748 8634 6776 9318
rect 6840 8906 6868 9646
rect 7104 9590 7156 9596
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6932 9042 6960 9386
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 7116 8786 7144 9590
rect 7208 9178 7236 10542
rect 7300 10266 7328 10542
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6840 8758 7144 8786
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6644 7200 6696 7206
rect 6564 7160 6644 7188
rect 6644 7142 6696 7148
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6564 5624 6592 6938
rect 6656 5846 6684 7142
rect 6748 5914 6776 8434
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5840 6696 5846
rect 6840 5794 6868 8758
rect 7208 8634 7236 9114
rect 7300 8974 7328 9998
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7392 8566 7420 11290
rect 7760 11286 7788 11494
rect 7748 11280 7800 11286
rect 7668 11240 7748 11268
rect 7668 10742 7696 11240
rect 7748 11222 7800 11228
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 8220 9908 8248 15098
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8312 13530 8340 14350
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13394 8432 14214
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8496 13326 8524 14214
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8588 13530 8616 14010
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8680 13258 8708 13806
rect 8772 13530 8800 16526
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12102 8340 12718
rect 8404 12714 8432 13194
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8588 12753 8616 12922
rect 8574 12744 8630 12753
rect 8392 12708 8444 12714
rect 8574 12679 8630 12688
rect 8392 12650 8444 12656
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8484 12232 8536 12238
rect 8404 12180 8484 12186
rect 8404 12174 8536 12180
rect 8404 12158 8524 12174
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11898 8340 12038
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8404 11830 8432 12158
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11898 8524 12038
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 7484 9880 8248 9908
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 6338 6960 7958
rect 7024 7002 7052 8366
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7116 7818 7144 8026
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7300 7478 7328 7822
rect 7392 7478 7420 7822
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7116 6934 7144 7142
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6390 7236 6598
rect 7392 6458 7420 7414
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7196 6384 7248 6390
rect 6932 6310 7052 6338
rect 7196 6326 7248 6332
rect 7024 6254 7052 6310
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6644 5782 6696 5788
rect 6748 5766 6868 5794
rect 6564 5596 6684 5624
rect 6656 5370 6684 5596
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6550 4992 6606 5001
rect 6550 4927 6606 4936
rect 6564 4457 6592 4927
rect 6550 4448 6606 4457
rect 6550 4383 6606 4392
rect 5908 4140 5960 4146
rect 6472 4134 6684 4162
rect 5908 4082 5960 4088
rect 6552 4072 6604 4078
rect 5998 4040 6054 4049
rect 6552 4014 6604 4020
rect 5998 3975 6054 3984
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5644 3182 5764 3210
rect 5540 2984 5592 2990
rect 5592 2944 5672 2972
rect 5540 2926 5592 2932
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2650 5580 2790
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5552 2514 5580 2586
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5644 2446 5672 2944
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 4908 2038 4936 2382
rect 5276 2310 5304 2382
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 4896 2032 4948 2038
rect 4896 1974 4948 1980
rect 4804 1896 4856 1902
rect 5368 1873 5396 2382
rect 4804 1838 4856 1844
rect 5354 1864 5410 1873
rect 5354 1799 5410 1808
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5000 800 5028 1294
rect 5736 800 5764 3182
rect 2686 776 2742 785
rect 2686 711 2742 720
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6012 762 6040 3975
rect 6276 3936 6328 3942
rect 6328 3896 6500 3924
rect 6276 3878 6328 3884
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 6472 2446 6500 3896
rect 6564 3505 6592 4014
rect 6656 3738 6684 4134
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6550 3496 6606 3505
rect 6550 3431 6606 3440
rect 6564 3194 6592 3431
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6656 3058 6684 3674
rect 6748 3058 6776 5766
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5370 6868 5646
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6932 5234 6960 6190
rect 7102 6080 7158 6089
rect 7102 6015 7158 6024
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6840 5137 6868 5170
rect 6826 5128 6882 5137
rect 7024 5114 7052 5646
rect 7116 5234 7144 6015
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7208 5794 7236 5850
rect 7392 5846 7420 6258
rect 7484 5914 7512 9880
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7748 9580 7800 9586
rect 7576 9540 7748 9568
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7380 5840 7432 5846
rect 7208 5766 7328 5794
rect 7380 5782 7432 5788
rect 7196 5704 7248 5710
rect 7300 5692 7328 5766
rect 7300 5664 7420 5692
rect 7196 5646 7248 5652
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7024 5086 7144 5114
rect 6826 5063 6882 5072
rect 6918 4856 6974 4865
rect 6828 4820 6880 4826
rect 6918 4791 6974 4800
rect 6828 4762 6880 4768
rect 6840 4214 6868 4762
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6932 3126 6960 4791
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7024 4282 7052 4490
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 3584 7052 4082
rect 7116 4078 7144 5086
rect 7208 4078 7236 5646
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7300 3942 7328 4422
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7116 3738 7144 3878
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7024 3556 7144 3584
rect 7116 3466 7144 3556
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7024 3194 7052 3402
rect 7208 3194 7236 3878
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 7392 2990 7420 5664
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3670 7512 3878
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7196 2984 7248 2990
rect 7024 2932 7196 2938
rect 7024 2926 7248 2932
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7024 2922 7236 2926
rect 7012 2916 7236 2922
rect 7064 2910 7236 2916
rect 7012 2858 7064 2864
rect 6642 2680 6698 2689
rect 6642 2615 6698 2624
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6656 2310 6684 2615
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 2106 6776 2246
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 7116 1601 7144 2314
rect 7208 1834 7236 2314
rect 7196 1828 7248 1834
rect 7196 1770 7248 1776
rect 7102 1592 7158 1601
rect 7102 1527 7158 1536
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 7208 870 7328 898
rect 7208 800 7236 870
rect 6012 734 6408 762
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7300 762 7328 870
rect 7576 762 7604 9540
rect 7748 9522 7800 9528
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7668 9178 7696 9386
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7944 8945 7972 9318
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 7930 8936 7986 8945
rect 7930 8871 7986 8880
rect 7748 8832 7800 8838
rect 7668 8792 7748 8820
rect 7668 7886 7696 8792
rect 7748 8774 7800 8780
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 6730 7696 7686
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 8220 7478 8248 8230
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7760 5710 7788 6394
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5914 7880 6190
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5704 7800 5710
rect 8220 5681 8248 7414
rect 8312 7342 8340 8434
rect 8404 7970 8432 11766
rect 8484 11144 8536 11150
rect 8482 11112 8484 11121
rect 8536 11112 8538 11121
rect 8482 11047 8538 11056
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10674 8524 10950
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8680 9466 8708 12582
rect 8772 10742 8800 13466
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9048 12238 9076 12650
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8956 11354 8984 12174
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10810 8892 11086
rect 8956 10810 8984 11290
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 9048 9654 9076 9959
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 9140 9518 9168 14758
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9876 14550 9904 16594
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9968 15094 9996 16050
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9324 13818 9352 14282
rect 9508 14074 9536 14282
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9876 13870 9904 14486
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 13864 9916 13870
rect 9232 12850 9260 13806
rect 9324 13790 9444 13818
rect 9864 13806 9916 13812
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9324 13258 9352 13670
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 12442 9260 12786
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9416 10810 9444 13790
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 9968 11014 9996 14418
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9220 10600 9272 10606
rect 9416 10554 9444 10746
rect 10060 10674 10088 12038
rect 10152 11762 10180 12582
rect 10244 12322 10272 14554
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10336 13530 10364 13874
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10244 12294 10364 12322
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10244 11898 10272 12174
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 10668 10100 10674
rect 9220 10542 9272 10548
rect 9232 10130 9260 10542
rect 9324 10526 9444 10554
rect 9876 10628 10048 10656
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9324 10062 9352 10526
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10266 9444 10406
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9404 10260 9456 10266
rect 9876 10248 9904 10628
rect 10048 10610 10100 10616
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9404 10202 9456 10208
rect 9508 10220 9904 10248
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9722 9444 9862
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9508 9568 9536 10220
rect 9772 10124 9824 10130
rect 9968 10112 9996 10406
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10060 10169 10088 10202
rect 9824 10084 9996 10112
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 9772 10066 9824 10072
rect 9680 10056 9732 10062
rect 10336 10010 10364 12294
rect 10428 11830 10456 12786
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10428 11200 10456 11766
rect 10796 11200 10824 14962
rect 10980 14414 11008 17138
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14646 16960 14702 16969
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 14074 11008 14350
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 11778 10916 13738
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11702 13288 11758 13297
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 11898 11008 12174
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10888 11750 11008 11778
rect 10428 11172 10548 11200
rect 10796 11172 10916 11200
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 10554 10456 11018
rect 10520 10674 10548 11172
rect 10692 11008 10744 11014
rect 10888 10996 10916 11172
rect 10692 10950 10744 10956
rect 10796 10968 10916 10996
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10428 10526 10548 10554
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10130 10456 10406
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 9680 9998 9732 10004
rect 9692 9874 9720 9998
rect 9772 9988 9824 9994
rect 10244 9982 10364 10010
rect 9824 9948 9904 9976
rect 9772 9930 9824 9936
rect 9876 9874 9904 9948
rect 9954 9888 10010 9897
rect 9692 9846 9812 9874
rect 9876 9846 9954 9874
rect 9784 9738 9812 9846
rect 9954 9823 10010 9832
rect 9784 9710 10180 9738
rect 9784 9586 9812 9710
rect 9954 9616 10010 9625
rect 9416 9540 9536 9568
rect 9772 9580 9824 9586
rect 9128 9512 9180 9518
rect 8576 9444 8628 9450
rect 8680 9438 9076 9466
rect 9128 9454 9180 9460
rect 8576 9386 8628 9392
rect 8588 8090 8616 9386
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 8906 8708 9318
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8850 8256 8906 8265
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8404 7942 8708 7970
rect 8574 7848 8630 7857
rect 8484 7812 8536 7818
rect 8574 7783 8630 7792
rect 8484 7754 8536 7760
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6118 8340 7142
rect 8404 6798 8432 7278
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8404 5710 8432 6734
rect 8496 6458 8524 7754
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8588 6338 8616 7783
rect 8496 6310 8616 6338
rect 8392 5704 8444 5710
rect 7748 5646 7800 5652
rect 8206 5672 8262 5681
rect 8392 5646 8444 5652
rect 8206 5607 8262 5616
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 4010 7696 5510
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 8220 5302 8248 5607
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8404 5098 8432 5646
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 8312 4282 8340 4966
rect 8404 4690 8432 5034
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8404 4282 8432 4490
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8496 4078 8524 6310
rect 8574 5128 8630 5137
rect 8574 5063 8630 5072
rect 8588 4690 8616 5063
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 7748 4072 7800 4078
rect 8484 4072 8536 4078
rect 7748 4014 7800 4020
rect 8390 4040 8446 4049
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7760 3738 7788 4014
rect 8484 4014 8536 4020
rect 8390 3975 8446 3984
rect 8576 4004 8628 4010
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7852 3398 7880 3674
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7654 3224 7710 3233
rect 7803 3227 8111 3236
rect 7654 3159 7710 3168
rect 7668 3126 7696 3159
rect 8220 3126 8248 3538
rect 7656 3120 7708 3126
rect 8208 3120 8260 3126
rect 7656 3062 7708 3068
rect 7930 3088 7986 3097
rect 7668 2514 7696 3062
rect 8208 3062 8260 3068
rect 8312 3058 8340 3538
rect 8404 3369 8432 3975
rect 8576 3946 8628 3952
rect 8588 3466 8616 3946
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8390 3360 8446 3369
rect 8390 3295 8446 3304
rect 7930 3023 7932 3032
rect 7984 3023 7986 3032
rect 8300 3052 8352 3058
rect 7932 2994 7984 3000
rect 8300 2994 8352 3000
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7932 2848 7984 2854
rect 7746 2816 7802 2825
rect 7932 2790 7984 2796
rect 7746 2751 7802 2760
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7760 2360 7788 2751
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7852 2446 7880 2586
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7300 734 7604 762
rect 7668 2332 7788 2360
rect 7944 2360 7972 2790
rect 8128 2514 8156 2926
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7944 2332 8248 2360
rect 7668 762 7696 2332
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 8220 1766 8248 2332
rect 8312 2038 8340 2994
rect 8680 2774 8708 7942
rect 8772 7750 8800 8230
rect 8850 8191 8906 8200
rect 8864 8090 8892 8191
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8956 7970 8984 8298
rect 8864 7942 8984 7970
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6322 8800 6598
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8864 6089 8892 7942
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7002 8984 7822
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9048 6712 9076 9438
rect 9140 7886 9168 9454
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7954 9260 8230
rect 9324 8090 9352 9386
rect 9416 9024 9444 9540
rect 9954 9551 10010 9560
rect 9772 9522 9824 9528
rect 9496 9444 9548 9450
rect 9772 9444 9824 9450
rect 9548 9404 9772 9432
rect 9496 9386 9548 9392
rect 9772 9386 9824 9392
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9416 8996 9536 9024
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9310 7984 9366 7993
rect 9220 7948 9272 7954
rect 9310 7919 9366 7928
rect 9220 7890 9272 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9220 6724 9272 6730
rect 9048 6684 9220 6712
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6254 8984 6598
rect 9140 6322 9168 6684
rect 9220 6666 9272 6672
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8944 6248 8996 6254
rect 9324 6202 9352 7919
rect 9416 7868 9444 8842
rect 9508 8537 9536 8996
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9494 8528 9550 8537
rect 9494 8463 9550 8472
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 8294 9720 8434
rect 9680 8288 9732 8294
rect 9784 8276 9812 8774
rect 9968 8634 9996 9551
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9110 10088 9318
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10060 8514 10088 9046
rect 9876 8498 10088 8514
rect 9864 8492 10088 8498
rect 9916 8486 10088 8492
rect 9864 8434 9916 8440
rect 9784 8248 9904 8276
rect 9680 8230 9732 8236
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9588 7880 9640 7886
rect 9416 7840 9588 7868
rect 9588 7822 9640 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 8944 6190 8996 6196
rect 9140 6174 9352 6202
rect 8850 6080 8906 6089
rect 8850 6015 8906 6024
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 4434 8800 5782
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8772 4406 8892 4434
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8772 3126 8800 4218
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8864 2774 8892 4406
rect 8956 3602 8984 4558
rect 9048 4282 9076 4694
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9048 3194 9076 3878
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9140 2774 9168 6174
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9232 4706 9260 5034
rect 9416 4808 9444 7686
rect 9600 7546 9628 7822
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9508 6225 9536 6938
rect 9876 6458 9904 8248
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 7206 9996 7890
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9494 6216 9550 6225
rect 9494 6151 9550 6160
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 10060 5778 10088 7958
rect 10152 6254 10180 9710
rect 10244 7528 10272 9982
rect 10520 9654 10548 10526
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9897 10640 10134
rect 10598 9888 10654 9897
rect 10598 9823 10654 9832
rect 10508 9648 10560 9654
rect 10414 9616 10470 9625
rect 10508 9590 10560 9596
rect 10414 9551 10416 9560
rect 10468 9551 10470 9560
rect 10416 9522 10468 9528
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10336 8634 10364 9454
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 8634 10456 9386
rect 10508 9376 10560 9382
rect 10560 9336 10640 9364
rect 10508 9318 10560 9324
rect 10506 9208 10562 9217
rect 10506 9143 10562 9152
rect 10520 9042 10548 9143
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10612 8906 10640 9336
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8832 10560 8838
rect 10560 8780 10640 8786
rect 10508 8774 10640 8780
rect 10520 8758 10640 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10520 8362 10548 8502
rect 10612 8362 10640 8758
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10244 7500 10364 7528
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 6730 10272 7346
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10152 5846 10180 6190
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9876 4826 9904 5578
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9968 5114 9996 5306
rect 10060 5234 10272 5250
rect 10048 5228 10272 5234
rect 10100 5222 10272 5228
rect 10048 5170 10100 5176
rect 9968 5086 10180 5114
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9864 4820 9916 4826
rect 9416 4780 9536 4808
rect 9232 4678 9444 4706
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 4146 9260 4558
rect 9416 4146 9444 4678
rect 9508 4554 9536 4780
rect 9864 4762 9916 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9876 4593 9904 4626
rect 9862 4584 9918 4593
rect 9496 4548 9548 4554
rect 9862 4519 9918 4528
rect 9496 4490 9548 4496
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9232 3126 9260 4082
rect 9416 3534 9444 4082
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 8496 2746 8708 2774
rect 8772 2746 8892 2774
rect 8956 2746 9168 2774
rect 8496 2038 8524 2746
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8588 2378 8616 2518
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8300 2032 8352 2038
rect 8300 1974 8352 1980
rect 8484 2032 8536 2038
rect 8484 1974 8536 1980
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 7852 870 7972 898
rect 7852 762 7880 870
rect 7944 800 7972 870
rect 8680 800 8708 2246
rect 8772 2038 8800 2746
rect 8760 2032 8812 2038
rect 8760 1974 8812 1980
rect 8956 1698 8984 2746
rect 9232 2689 9260 2858
rect 9416 2854 9444 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9600 2990 9628 3130
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9218 2680 9274 2689
rect 9517 2683 9825 2692
rect 9218 2615 9274 2624
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9034 2544 9090 2553
rect 9034 2479 9090 2488
rect 9048 2446 9076 2479
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 8944 1692 8996 1698
rect 8944 1634 8996 1640
rect 9416 800 9444 2314
rect 9692 1714 9720 2586
rect 9770 2544 9826 2553
rect 9770 2479 9772 2488
rect 9824 2479 9826 2488
rect 9772 2450 9824 2456
rect 9876 2394 9904 4150
rect 9784 2366 9904 2394
rect 9784 1834 9812 2366
rect 9968 2038 9996 4966
rect 9956 2032 10008 2038
rect 9956 1974 10008 1980
rect 9772 1828 9824 1834
rect 9772 1770 9824 1776
rect 10060 1714 10088 4966
rect 10152 4282 10180 5086
rect 10244 4690 10272 5222
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10336 4321 10364 7500
rect 10612 7460 10640 8298
rect 10520 7432 10640 7460
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 5658 10456 6802
rect 10520 6186 10548 7432
rect 10704 6882 10732 10950
rect 10796 8634 10824 10968
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10980 10554 11008 11750
rect 11072 11150 11100 13262
rect 11702 13223 11758 13232
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11532 12306 11560 12854
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11164 11898 11192 12174
rect 11624 12170 11652 13126
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10674 11100 11086
rect 11716 10996 11744 13223
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 11121 11836 12922
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11900 11354 11928 11698
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11900 11218 11928 11290
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11794 11112 11850 11121
rect 11794 11047 11850 11056
rect 11716 10968 11836 10996
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11152 10600 11204 10606
rect 10888 10266 10916 10542
rect 10980 10526 11100 10554
rect 11152 10542 11204 10548
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10888 8537 10916 9522
rect 10980 9110 11008 9862
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11072 8922 11100 10526
rect 11164 9568 11192 10542
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10266 11376 10406
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 11244 9580 11296 9586
rect 11164 9540 11244 9568
rect 11244 9522 11296 9528
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10980 8894 11100 8922
rect 10874 8528 10930 8537
rect 10784 8492 10836 8498
rect 10874 8463 10930 8472
rect 10784 8434 10836 8440
rect 10796 8294 10824 8434
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10980 7313 11008 8894
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 7750 11100 8774
rect 11164 8362 11192 8978
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11624 8498 11652 10610
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9722 11744 9998
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11716 9178 11744 9454
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11702 8664 11758 8673
rect 11702 8599 11704 8608
rect 11756 8599 11758 8608
rect 11704 8570 11756 8576
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7857 11376 8230
rect 11624 7886 11652 8434
rect 11702 7984 11758 7993
rect 11702 7919 11758 7928
rect 11612 7880 11664 7886
rect 11334 7848 11390 7857
rect 11612 7822 11664 7828
rect 11334 7783 11390 7792
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10966 7304 11022 7313
rect 10966 7239 11022 7248
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10612 6854 10732 6882
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10428 5630 10548 5658
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10322 4312 10378 4321
rect 10140 4276 10192 4282
rect 10322 4247 10378 4256
rect 10140 4218 10192 4224
rect 10428 3754 10456 5510
rect 10336 3726 10456 3754
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9692 1686 10088 1714
rect 9954 1456 10010 1465
rect 9954 1391 10010 1400
rect 9968 1358 9996 1391
rect 9956 1352 10008 1358
rect 9956 1294 10008 1300
rect 10152 800 10180 2790
rect 10230 2544 10286 2553
rect 10336 2514 10364 3726
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10230 2479 10286 2488
rect 10324 2508 10376 2514
rect 10244 1290 10272 2479
rect 10324 2450 10376 2456
rect 10428 2446 10456 3606
rect 10520 2650 10548 5630
rect 10612 4826 10640 6854
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10980 6458 11008 7142
rect 11072 6644 11100 7686
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 11716 7392 11744 7919
rect 11624 7364 11744 7392
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6769 11192 7142
rect 11624 7002 11652 7364
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11150 6760 11206 6769
rect 11150 6695 11206 6704
rect 11072 6616 11192 6644
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10704 5137 10732 6122
rect 10980 5914 11008 6122
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5914 11100 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10968 5704 11020 5710
rect 10782 5672 10838 5681
rect 10968 5646 11020 5652
rect 10782 5607 10838 5616
rect 10690 5128 10746 5137
rect 10690 5063 10746 5072
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 4214 10640 4626
rect 10690 4584 10746 4593
rect 10690 4519 10746 4528
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10704 3754 10732 4519
rect 10612 3726 10732 3754
rect 10612 3670 10640 3726
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10704 3534 10732 3606
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10704 3058 10732 3470
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10796 2774 10824 5607
rect 10980 5370 11008 5646
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10980 4622 11008 4762
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11072 3777 11100 5034
rect 11058 3768 11114 3777
rect 11058 3703 11114 3712
rect 11164 3584 11192 6616
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5817 11284 6326
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5914 11468 6054
rect 11624 5914 11652 6802
rect 11716 6730 11744 7210
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6458 11744 6666
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11702 6352 11758 6361
rect 11702 6287 11704 6296
rect 11756 6287 11758 6296
rect 11704 6258 11756 6264
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11242 5808 11298 5817
rect 11242 5743 11298 5752
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11716 5234 11744 6122
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4826 11284 5102
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11072 3556 11192 3584
rect 10874 3360 10930 3369
rect 11072 3346 11100 3556
rect 11256 3448 11284 4082
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3618 11376 3878
rect 11440 3738 11468 4150
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11532 3618 11560 4014
rect 11624 3738 11652 5170
rect 11808 5114 11836 10968
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11992 9382 12020 9998
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11900 8974 11928 9318
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8634 11928 8774
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11900 7206 11928 8026
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11900 6254 11928 6802
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 5166 11928 6190
rect 11992 5778 12020 9318
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11992 5409 12020 5578
rect 11978 5400 12034 5409
rect 12084 5370 12112 15030
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 13740 14074 13768 16390
rect 13832 15706 13860 16390
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13394 12756 13670
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11150 12204 12242
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12176 10062 12204 10746
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9722 12204 9862
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12164 9512 12216 9518
rect 12162 9480 12164 9489
rect 12216 9480 12218 9489
rect 12162 9415 12218 9424
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 5794 12204 8230
rect 12268 6361 12296 13194
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12918 12664 13126
rect 13004 12986 13032 13262
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12306 12480 12582
rect 12728 12434 12756 12650
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 12544 12406 12756 12434
rect 12992 12436 13044 12442
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12360 9602 12388 12106
rect 12544 11200 12572 12406
rect 13280 12434 13308 12582
rect 13464 12442 13492 13126
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13452 12436 13504 12442
rect 13280 12406 13400 12434
rect 12992 12378 13044 12384
rect 13004 11694 13032 12378
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 11898 13216 12174
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12452 11172 12572 11200
rect 12452 9738 12480 11172
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10742 12664 10950
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12728 10554 12756 11562
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 13280 11354 13308 11698
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13372 11234 13400 12406
rect 13452 12378 13504 12384
rect 13280 11206 13400 11234
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12636 10526 12756 10554
rect 12636 9926 12664 10526
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 9994 12756 10406
rect 12820 10130 12848 10950
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13188 10577 13216 10678
rect 13174 10568 13230 10577
rect 13174 10503 13230 10512
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 13084 10056 13136 10062
rect 13176 10056 13228 10062
rect 13084 9998 13136 10004
rect 13174 10024 13176 10033
rect 13228 10024 13230 10033
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12452 9710 12572 9738
rect 12360 9574 12480 9602
rect 12452 7970 12480 9574
rect 12360 7942 12480 7970
rect 12360 7290 12388 7942
rect 12544 7426 12572 9710
rect 12728 9654 12756 9930
rect 12912 9722 12940 9930
rect 13096 9722 13124 9998
rect 13174 9959 13230 9968
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12636 9178 12664 9522
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12820 9058 12848 9522
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 12728 9030 12848 9058
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8634 12664 8774
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8514 12756 9030
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12636 8486 12756 8514
rect 12636 7750 12664 8486
rect 12820 7886 12848 8774
rect 12912 8634 12940 8910
rect 13280 8786 13308 11206
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13372 9654 13400 11018
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10198 13492 10542
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 9042 13400 9318
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13556 8922 13584 12582
rect 13924 12434 13952 15438
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13924 12406 14044 12434
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11898 13676 12038
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13648 11354 13676 11834
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10538 13676 10950
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13648 9926 13676 10474
rect 13740 10130 13768 11222
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 8968 13780 8974
rect 13556 8894 13676 8922
rect 13728 8910 13780 8916
rect 13452 8832 13504 8838
rect 13280 8758 13400 8786
rect 13452 8774 13504 8780
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12912 8498 12940 8570
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12544 7398 12664 7426
rect 12360 7262 12572 7290
rect 12254 6352 12310 6361
rect 12254 6287 12310 6296
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5914 12296 6054
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12176 5766 12296 5794
rect 11978 5335 12034 5344
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11716 5086 11836 5114
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11716 4078 11744 5086
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11348 3590 11560 3618
rect 11610 3632 11666 3641
rect 11348 3505 11376 3590
rect 11610 3567 11666 3576
rect 11624 3534 11652 3567
rect 11612 3528 11664 3534
rect 10874 3295 10930 3304
rect 10980 3318 11100 3346
rect 11164 3420 11284 3448
rect 11334 3496 11390 3505
rect 11612 3470 11664 3476
rect 11334 3431 11390 3440
rect 10888 2990 10916 3295
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10612 2746 10824 2774
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10232 1284 10284 1290
rect 10232 1226 10284 1232
rect 7668 734 7880 762
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10612 762 10640 2746
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10796 2514 10824 2615
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10980 2310 11008 3318
rect 11164 3176 11192 3420
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11244 3188 11296 3194
rect 11164 3148 11244 3176
rect 11244 3130 11296 3136
rect 11624 3058 11652 3470
rect 11716 3194 11744 3878
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11164 1970 11192 2382
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 11256 1465 11284 1702
rect 11242 1456 11298 1465
rect 11242 1391 11298 1400
rect 10796 870 10916 898
rect 10796 762 10824 870
rect 10888 800 10916 870
rect 11624 800 11652 2858
rect 11704 2372 11756 2378
rect 11808 2360 11836 4966
rect 11900 3602 11928 5102
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11992 4185 12020 4490
rect 11978 4176 12034 4185
rect 11978 4111 12034 4120
rect 12084 4078 12112 4626
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11992 3618 12020 4014
rect 12084 3738 12112 4014
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12162 3632 12218 3641
rect 11888 3596 11940 3602
rect 11992 3590 12112 3618
rect 11888 3538 11940 3544
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11900 3194 11928 3402
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11992 2582 12020 3402
rect 11980 2576 12032 2582
rect 11886 2544 11942 2553
rect 11980 2518 12032 2524
rect 11886 2479 11942 2488
rect 11900 2378 11928 2479
rect 12084 2417 12112 3590
rect 12162 3567 12218 3576
rect 12176 2990 12204 3567
rect 12268 3194 12296 5766
rect 12346 5672 12402 5681
rect 12346 5607 12348 5616
rect 12400 5607 12402 5616
rect 12348 5578 12400 5584
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 4826 12480 5510
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12360 3369 12388 4014
rect 12346 3360 12402 3369
rect 12346 3295 12402 3304
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12070 2408 12126 2417
rect 11756 2332 11836 2360
rect 11888 2372 11940 2378
rect 11704 2314 11756 2320
rect 12452 2378 12480 4762
rect 12544 3126 12572 7262
rect 12636 6730 12664 7398
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12622 6488 12678 6497
rect 12622 6423 12678 6432
rect 12636 5710 12664 6423
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12728 5302 12756 7754
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7342 12848 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12820 6390 12848 7278
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 13280 6798 13308 7142
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 13096 6254 13124 6666
rect 13372 6610 13400 8758
rect 13464 7818 13492 8774
rect 13556 8673 13584 8774
rect 13542 8664 13598 8673
rect 13542 8599 13598 8608
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13556 7818 13584 8298
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13280 6582 13400 6610
rect 13084 6248 13136 6254
rect 12820 6196 13084 6202
rect 12820 6190 13136 6196
rect 12820 6174 13124 6190
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12636 3942 12664 5238
rect 12820 4690 12848 6174
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 13280 4706 13308 6582
rect 13464 5914 13492 7414
rect 13556 6934 13584 7754
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13556 6458 13584 6734
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13648 5302 13676 8894
rect 13740 7177 13768 8910
rect 13832 8498 13860 9318
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13726 7168 13782 7177
rect 13726 7103 13782 7112
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13372 4826 13400 5170
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 12808 4684 12860 4690
rect 13280 4678 13400 4706
rect 12808 4626 12860 4632
rect 13096 4146 13216 4162
rect 13372 4146 13400 4678
rect 13464 4593 13492 4966
rect 13740 4826 13768 6870
rect 13832 6866 13860 7890
rect 13924 7886 13952 8366
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 7546 13952 7822
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6254 13860 6598
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13924 5846 13952 7142
rect 14016 6798 14044 12406
rect 14108 10470 14136 13874
rect 14292 13530 14320 16934
rect 14646 16895 14702 16904
rect 14660 16794 14688 16895
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 15028 16153 15056 16526
rect 15014 16144 15070 16153
rect 15014 16079 15070 16088
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14844 15473 14872 15574
rect 14830 15464 14886 15473
rect 14830 15399 14886 15408
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14521 14412 14758
rect 14370 14512 14426 14521
rect 14370 14447 14426 14456
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13705 14504 13806
rect 14462 13696 14518 13705
rect 14462 13631 14518 13640
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14200 12442 14228 13262
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12889 14412 13126
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14188 12232 14240 12238
rect 14384 12209 14412 12310
rect 14188 12174 14240 12180
rect 14370 12200 14426 12209
rect 14200 11898 14228 12174
rect 14370 12135 14426 12144
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14292 11150 14320 11494
rect 14384 11257 14412 11494
rect 14370 11248 14426 11257
rect 14370 11183 14426 11192
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14186 10568 14242 10577
rect 14186 10503 14242 10512
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14200 9722 14228 10503
rect 14370 10432 14426 10441
rect 14370 10367 14426 10376
rect 14384 10266 14412 10367
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14476 10146 14504 12718
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14292 10118 14504 10146
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14094 9616 14150 9625
rect 14094 9551 14096 9560
rect 14148 9551 14150 9560
rect 14096 9522 14148 9528
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8090 14136 9046
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13726 4720 13782 4729
rect 13726 4655 13782 4664
rect 13636 4616 13688 4622
rect 13450 4584 13506 4593
rect 13636 4558 13688 4564
rect 13450 4519 13506 4528
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13084 4140 13216 4146
rect 13136 4134 13216 4140
rect 13084 4082 13136 4088
rect 13188 4026 13216 4134
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13188 3998 13308 4026
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12716 2984 12768 2990
rect 12530 2952 12586 2961
rect 12716 2926 12768 2932
rect 12530 2887 12586 2896
rect 12544 2378 12572 2887
rect 12070 2343 12126 2352
rect 12440 2372 12492 2378
rect 11888 2314 11940 2320
rect 12440 2314 12492 2320
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12176 2038 12204 2246
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12728 1902 12756 2926
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12820 2514 12848 2586
rect 13280 2514 13308 3998
rect 13464 3534 13492 4422
rect 13556 4282 13584 4490
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13648 3194 13676 4558
rect 13740 3534 13768 4655
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13372 2582 13400 3062
rect 13832 2922 13860 4422
rect 13924 4146 13952 5782
rect 14016 4214 14044 6054
rect 14108 5370 14136 7142
rect 14200 5370 14228 8366
rect 14292 7002 14320 10118
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14384 8945 14412 9046
rect 14370 8936 14426 8945
rect 14370 8871 14426 8880
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 6458 14412 8502
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14200 4060 14228 4966
rect 14108 4032 14228 4060
rect 14108 3738 14136 4032
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12348 1284 12400 1290
rect 12348 1226 12400 1232
rect 12360 800 12388 1226
rect 13096 800 13124 2042
rect 13832 870 13952 898
rect 13832 800 13860 870
rect 10612 734 10824 762
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 13924 762 13952 870
rect 14200 762 14228 3878
rect 14292 2650 14320 5646
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14384 5098 14412 5578
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 3602 14412 5034
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14476 3482 14504 9998
rect 14568 5574 14596 12582
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14384 3454 14504 3482
rect 14556 3460 14608 3466
rect 14384 2990 14412 3454
rect 14556 3402 14608 3408
rect 14462 3088 14518 3097
rect 14462 3023 14464 3032
rect 14516 3023 14518 3032
rect 14464 2994 14516 3000
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14278 2544 14334 2553
rect 14278 2479 14334 2488
rect 14292 2446 14320 2479
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 14568 800 14596 3402
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 13924 734 14228 762
rect 14554 0 14610 800
<< via2 >>
rect 2778 18536 2834 18592
rect 13726 18536 13782 18592
rect 938 17720 994 17776
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 14646 17720 14702 17776
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 1030 16940 1032 16960
rect 1032 16940 1084 16960
rect 1084 16940 1086 16960
rect 1030 16904 1086 16940
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 938 16088 994 16144
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 1122 15272 1178 15328
rect 1582 14592 1638 14648
rect 1490 14320 1546 14376
rect 570 3304 626 3360
rect 938 12824 994 12880
rect 1030 12280 1086 12336
rect 938 12044 940 12064
rect 940 12044 992 12064
rect 992 12044 994 12064
rect 938 12008 994 12044
rect 938 10376 994 10432
rect 938 9560 994 9616
rect 938 4664 994 4720
rect 1582 13676 1584 13696
rect 1584 13676 1636 13696
rect 1636 13676 1638 13696
rect 1582 13640 1638 13676
rect 1582 12588 1584 12608
rect 1584 12588 1636 12608
rect 1636 12588 1638 12608
rect 1582 12552 1638 12588
rect 1674 11092 1676 11112
rect 1676 11092 1728 11112
rect 1728 11092 1730 11112
rect 1674 11056 1730 11092
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2410 14476 2466 14512
rect 2410 14456 2412 14476
rect 2412 14456 2464 14476
rect 2464 14456 2466 14476
rect 2318 13776 2374 13832
rect 2042 11600 2098 11656
rect 1858 10648 1914 10704
rect 1490 7928 1546 7984
rect 1490 7812 1546 7848
rect 1490 7792 1492 7812
rect 1492 7792 1544 7812
rect 1544 7792 1546 7812
rect 1490 7248 1546 7304
rect 1398 6296 1454 6352
rect 1306 5208 1362 5264
rect 1858 8336 1914 8392
rect 1674 5480 1730 5536
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 2962 12708 3018 12744
rect 2962 12688 2964 12708
rect 2964 12688 3016 12708
rect 3016 12688 3018 12708
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 3238 14184 3294 14240
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 3238 13232 3294 13288
rect 3330 12960 3386 13016
rect 3238 12588 3240 12608
rect 3240 12588 3292 12608
rect 3292 12588 3294 12608
rect 3238 12552 3294 12588
rect 3054 12008 3110 12064
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 3054 11056 3110 11112
rect 2318 10784 2374 10840
rect 2318 10512 2374 10568
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 2318 9424 2374 9480
rect 2226 9016 2282 9072
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 2042 6840 2098 6896
rect 2318 7928 2374 7984
rect 2594 8336 2650 8392
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 1950 4528 2006 4584
rect 1490 2916 1546 2952
rect 1490 2896 1492 2916
rect 1492 2896 1544 2916
rect 1544 2896 1546 2916
rect 2226 4120 2282 4176
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 2410 4020 2412 4040
rect 2412 4020 2464 4040
rect 2464 4020 2466 4040
rect 2410 3984 2466 4020
rect 2962 3984 3018 4040
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 3422 9868 3424 9888
rect 3424 9868 3476 9888
rect 3476 9868 3478 9888
rect 3422 9832 3478 9868
rect 3422 9288 3478 9344
rect 4066 13776 4122 13832
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 4710 13776 4766 13832
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 3882 12552 3938 12608
rect 3790 12144 3846 12200
rect 3790 10784 3846 10840
rect 4066 11192 4122 11248
rect 4066 10648 4122 10704
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 4250 11600 4306 11656
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4710 9016 4766 9072
rect 3974 7656 4030 7712
rect 3882 6976 3938 7032
rect 3974 6024 4030 6080
rect 3330 3848 3386 3904
rect 3238 3440 3294 3496
rect 3238 3304 3294 3360
rect 3514 5072 3570 5128
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 4710 8472 4766 8528
rect 4434 8064 4490 8120
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 4986 12960 5042 13016
rect 5262 13096 5318 13152
rect 5170 12824 5226 12880
rect 4894 10240 4950 10296
rect 4618 6296 4674 6352
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 3790 3712 3846 3768
rect 3882 3576 3938 3632
rect 3882 3440 3938 3496
rect 3146 2624 3202 2680
rect 2594 2488 2650 2544
rect 3330 2352 3386 2408
rect 4066 4120 4122 4176
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 5170 12280 5226 12336
rect 5262 11736 5318 11792
rect 5078 7384 5134 7440
rect 5538 12688 5594 12744
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 5814 12724 5816 12744
rect 5816 12724 5868 12744
rect 5868 12724 5870 12744
rect 5814 12688 5870 12724
rect 5722 12552 5778 12608
rect 5630 10240 5686 10296
rect 5170 6024 5226 6080
rect 5078 5208 5134 5264
rect 4894 4392 4950 4448
rect 4802 4020 4804 4040
rect 4804 4020 4856 4040
rect 4856 4020 4858 4040
rect 4802 3984 4858 4020
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 4986 3052 5042 3088
rect 4986 3032 4988 3052
rect 4988 3032 5040 3052
rect 5040 3032 5042 3052
rect 4250 2760 4306 2816
rect 4066 2488 4122 2544
rect 5446 7928 5502 7984
rect 5630 9288 5686 9344
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6550 10104 6606 10160
rect 6918 11736 6974 11792
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 7102 11192 7158 11248
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 5906 8064 5962 8120
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 5814 5616 5870 5672
rect 5354 4664 5410 4720
rect 5262 3848 5318 3904
rect 4618 2624 4674 2680
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 6366 5752 6422 5808
rect 6182 5344 6238 5400
rect 6090 5072 6146 5128
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 5722 4256 5778 4312
rect 5722 3712 5778 3768
rect 5630 3576 5686 3632
rect 6366 4276 6422 4312
rect 6366 4256 6368 4276
rect 6368 4256 6420 4276
rect 6420 4256 6422 4276
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 8574 12688 8630 12744
rect 6550 4936 6606 4992
rect 6550 4392 6606 4448
rect 5998 3984 6054 4040
rect 5722 3304 5778 3360
rect 5354 1808 5410 1864
rect 2686 720 2742 776
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 6550 3440 6606 3496
rect 7102 6024 7158 6080
rect 6826 5072 6882 5128
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 6918 4800 6974 4856
rect 6642 2624 6698 2680
rect 7102 1536 7158 1592
rect 7930 8880 7986 8936
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 8482 11092 8484 11112
rect 8484 11092 8536 11112
rect 8536 11092 8538 11112
rect 8482 11056 8538 11092
rect 9034 9968 9090 10024
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 10046 10104 10102 10160
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 9954 9832 10010 9888
rect 8574 7792 8630 7848
rect 8206 5616 8262 5672
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 8574 5072 8630 5128
rect 8390 3984 8446 4040
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 7654 3168 7710 3224
rect 7930 3052 7986 3088
rect 8390 3304 8446 3360
rect 7930 3032 7932 3052
rect 7932 3032 7984 3052
rect 7984 3032 7986 3052
rect 7746 2760 7802 2816
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 8850 8200 8906 8256
rect 9954 9560 10010 9616
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 9310 7928 9366 7984
rect 9494 8472 9550 8528
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 8850 6024 8906 6080
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9494 6160 9550 6216
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 10598 9832 10654 9888
rect 10414 9580 10470 9616
rect 10414 9560 10416 9580
rect 10416 9560 10468 9580
rect 10468 9560 10470 9580
rect 10506 9152 10562 9208
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9862 4528 9918 4584
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 9218 2624 9274 2680
rect 9034 2488 9090 2544
rect 9770 2508 9826 2544
rect 9770 2488 9772 2508
rect 9772 2488 9824 2508
rect 9824 2488 9826 2508
rect 11702 13232 11758 13288
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 11794 11056 11850 11112
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 10874 8472 10930 8528
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11702 8628 11758 8664
rect 11702 8608 11704 8628
rect 11704 8608 11756 8628
rect 11756 8608 11758 8628
rect 11702 7928 11758 7984
rect 11334 7792 11390 7848
rect 10966 7248 11022 7304
rect 10322 4256 10378 4312
rect 9954 1400 10010 1456
rect 10230 2488 10286 2544
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 11150 6704 11206 6760
rect 10782 5616 10838 5672
rect 10690 5072 10746 5128
rect 10690 4528 10746 4584
rect 11058 3712 11114 3768
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11702 6316 11758 6352
rect 11702 6296 11704 6316
rect 11704 6296 11756 6316
rect 11756 6296 11758 6316
rect 11242 5752 11298 5808
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 10874 3304 10930 3360
rect 11978 5344 12034 5400
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 12162 9460 12164 9480
rect 12164 9460 12216 9480
rect 12216 9460 12218 9480
rect 12162 9424 12218 9460
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 13174 10512 13230 10568
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 13174 10004 13176 10024
rect 13176 10004 13228 10024
rect 13228 10004 13230 10024
rect 13174 9968 13230 10004
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 12254 6296 12310 6352
rect 11610 3576 11666 3632
rect 11334 3440 11390 3496
rect 10782 2624 10838 2680
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 11242 1400 11298 1456
rect 11978 4120 12034 4176
rect 11886 2488 11942 2544
rect 12162 3576 12218 3632
rect 12346 5636 12402 5672
rect 12346 5616 12348 5636
rect 12348 5616 12400 5636
rect 12400 5616 12402 5636
rect 12346 3304 12402 3360
rect 12070 2352 12126 2408
rect 12622 6432 12678 6488
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 13542 8608 13598 8664
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 13726 7112 13782 7168
rect 14646 16904 14702 16960
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 15014 16088 15070 16144
rect 14830 15408 14886 15464
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14370 14456 14426 14512
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14462 13640 14518 13696
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14370 12824 14426 12880
rect 14370 12144 14426 12200
rect 14370 11192 14426 11248
rect 14186 10512 14242 10568
rect 14370 10376 14426 10432
rect 14094 9580 14150 9616
rect 14094 9560 14096 9580
rect 14096 9560 14148 9580
rect 14148 9560 14150 9580
rect 13726 4664 13782 4720
rect 13450 4528 13506 4584
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 12530 2896 12586 2952
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14370 8880 14426 8936
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14462 3052 14518 3088
rect 14462 3032 14464 3052
rect 14464 3032 14516 3052
rect 14516 3032 14518 3052
rect 14278 2488 14334 2544
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
<< metal3 >>
rect 0 18594 800 18624
rect 2773 18594 2839 18597
rect 0 18592 2839 18594
rect 0 18536 2778 18592
rect 2834 18536 2839 18592
rect 0 18534 2839 18536
rect 0 18504 800 18534
rect 2773 18531 2839 18534
rect 13721 18594 13787 18597
rect 15200 18594 16000 18624
rect 13721 18592 16000 18594
rect 13721 18536 13726 18592
rect 13782 18536 16000 18592
rect 13721 18534 16000 18536
rect 13721 18531 13787 18534
rect 15200 18504 16000 18534
rect 0 17778 800 17808
rect 933 17778 999 17781
rect 0 17776 999 17778
rect 0 17720 938 17776
rect 994 17720 999 17776
rect 0 17718 999 17720
rect 0 17688 800 17718
rect 933 17715 999 17718
rect 14641 17778 14707 17781
rect 15200 17778 16000 17808
rect 14641 17776 16000 17778
rect 14641 17720 14646 17776
rect 14702 17720 16000 17776
rect 14641 17718 16000 17720
rect 14641 17715 14707 17718
rect 15200 17688 16000 17718
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 0 16962 800 16992
rect 1025 16962 1091 16965
rect 0 16960 1091 16962
rect 0 16904 1030 16960
rect 1086 16904 1091 16960
rect 0 16902 1091 16904
rect 0 16872 800 16902
rect 1025 16899 1091 16902
rect 14641 16962 14707 16965
rect 15200 16962 16000 16992
rect 14641 16960 16000 16962
rect 14641 16904 14646 16960
rect 14702 16904 16000 16960
rect 14641 16902 16000 16904
rect 14641 16899 14707 16902
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 15200 16872 16000 16902
rect 12940 16831 13256 16832
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 14653 16287 14969 16288
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 15009 16146 15075 16149
rect 15200 16146 16000 16176
rect 15009 16144 16000 16146
rect 15009 16088 15014 16144
rect 15070 16088 16000 16144
rect 15009 16086 16000 16088
rect 15009 16083 15075 16086
rect 15200 16056 16000 16086
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 14825 15466 14891 15469
rect 14825 15464 15210 15466
rect 14825 15408 14830 15464
rect 14886 15408 15210 15464
rect 14825 15406 15210 15408
rect 14825 15403 14891 15406
rect 15150 15360 15210 15406
rect 0 15330 800 15360
rect 1117 15330 1183 15333
rect 0 15328 1183 15330
rect 0 15272 1122 15328
rect 1178 15272 1183 15328
rect 0 15270 1183 15272
rect 15150 15270 16000 15360
rect 0 15240 800 15270
rect 1117 15267 1183 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 15200 15240 16000 15270
rect 14653 15199 14969 15200
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 1577 14650 1643 14653
rect 936 14648 1643 14650
rect 936 14592 1582 14648
rect 1638 14592 1643 14648
rect 936 14590 1643 14592
rect 0 14514 800 14544
rect 936 14514 996 14590
rect 1577 14587 1643 14590
rect 0 14454 996 14514
rect 2405 14514 2471 14517
rect 8334 14514 8340 14516
rect 2405 14512 8340 14514
rect 2405 14456 2410 14512
rect 2466 14456 8340 14512
rect 2405 14454 8340 14456
rect 0 14424 800 14454
rect 2405 14451 2471 14454
rect 8334 14452 8340 14454
rect 8404 14452 8410 14516
rect 14365 14514 14431 14517
rect 15200 14514 16000 14544
rect 14365 14512 16000 14514
rect 14365 14456 14370 14512
rect 14426 14456 16000 14512
rect 14365 14454 16000 14456
rect 14365 14451 14431 14454
rect 15200 14424 16000 14454
rect 1485 14378 1551 14381
rect 8518 14378 8524 14380
rect 1485 14376 8524 14378
rect 1485 14320 1490 14376
rect 1546 14320 8524 14376
rect 1485 14318 8524 14320
rect 1485 14315 1551 14318
rect 8518 14316 8524 14318
rect 8588 14316 8594 14380
rect 1158 14180 1164 14244
rect 1228 14242 1234 14244
rect 3233 14242 3299 14245
rect 1228 14240 3299 14242
rect 1228 14184 3238 14240
rect 3294 14184 3299 14240
rect 1228 14182 3299 14184
rect 1228 14180 1234 14182
rect 3233 14179 3299 14182
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 9070 13970 9076 13972
rect 4478 13910 9076 13970
rect 974 13772 980 13836
rect 1044 13834 1050 13836
rect 2313 13834 2379 13837
rect 1044 13832 2379 13834
rect 1044 13776 2318 13832
rect 2374 13776 2379 13832
rect 1044 13774 2379 13776
rect 1044 13772 1050 13774
rect 2313 13771 2379 13774
rect 4061 13834 4127 13837
rect 4478 13834 4538 13910
rect 9070 13908 9076 13910
rect 9140 13908 9146 13972
rect 4061 13832 4538 13834
rect 4061 13776 4066 13832
rect 4122 13776 4538 13832
rect 4061 13774 4538 13776
rect 4705 13834 4771 13837
rect 9990 13834 9996 13836
rect 4705 13832 9996 13834
rect 4705 13776 4710 13832
rect 4766 13776 9996 13832
rect 4705 13774 9996 13776
rect 4061 13771 4127 13774
rect 4705 13771 4771 13774
rect 9990 13772 9996 13774
rect 10060 13772 10066 13836
rect 0 13698 800 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 800 13638
rect 1577 13635 1643 13638
rect 14457 13698 14523 13701
rect 15200 13698 16000 13728
rect 14457 13696 16000 13698
rect 14457 13640 14462 13696
rect 14518 13640 16000 13696
rect 14457 13638 16000 13640
rect 14457 13635 14523 13638
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 15200 13608 16000 13638
rect 12940 13567 13256 13568
rect 3233 13290 3299 13293
rect 11697 13290 11763 13293
rect 3233 13288 11763 13290
rect 3233 13232 3238 13288
rect 3294 13232 11702 13288
rect 11758 13232 11763 13288
rect 3233 13230 11763 13232
rect 3233 13227 3299 13230
rect 11697 13227 11763 13230
rect 5257 13154 5323 13157
rect 6494 13154 6500 13156
rect 5257 13152 6500 13154
rect 5257 13096 5262 13152
rect 5318 13096 6500 13152
rect 5257 13094 6500 13096
rect 5257 13091 5323 13094
rect 6494 13092 6500 13094
rect 6564 13092 6570 13156
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 14653 13023 14969 13024
rect 3325 13018 3391 13021
rect 4102 13018 4108 13020
rect 3325 13016 4108 13018
rect 3325 12960 3330 13016
rect 3386 12960 4108 13016
rect 3325 12958 4108 12960
rect 3325 12955 3391 12958
rect 4102 12956 4108 12958
rect 4172 12956 4178 13020
rect 4981 13018 5047 13021
rect 5574 13018 5580 13020
rect 4981 13016 5580 13018
rect 4981 12960 4986 13016
rect 5042 12960 5580 13016
rect 4981 12958 5580 12960
rect 4981 12955 5047 12958
rect 5574 12956 5580 12958
rect 5644 12956 5650 13020
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 5165 12882 5231 12885
rect 7414 12882 7420 12884
rect 5165 12880 7420 12882
rect 5165 12824 5170 12880
rect 5226 12824 7420 12880
rect 5165 12822 7420 12824
rect 5165 12819 5231 12822
rect 7414 12820 7420 12822
rect 7484 12820 7490 12884
rect 14365 12882 14431 12885
rect 15200 12882 16000 12912
rect 14365 12880 16000 12882
rect 14365 12824 14370 12880
rect 14426 12824 16000 12880
rect 14365 12822 16000 12824
rect 14365 12819 14431 12822
rect 15200 12792 16000 12822
rect 2957 12746 3023 12749
rect 5533 12746 5599 12749
rect 2957 12744 5599 12746
rect 2957 12688 2962 12744
rect 3018 12688 5538 12744
rect 5594 12688 5599 12744
rect 2957 12686 5599 12688
rect 2957 12683 3023 12686
rect 5533 12683 5599 12686
rect 5809 12746 5875 12749
rect 8569 12746 8635 12749
rect 5809 12744 8635 12746
rect 5809 12688 5814 12744
rect 5870 12688 8574 12744
rect 8630 12688 8635 12744
rect 5809 12686 8635 12688
rect 5809 12683 5875 12686
rect 8569 12683 8635 12686
rect 1577 12610 1643 12613
rect 2078 12610 2084 12612
rect 1577 12608 2084 12610
rect 1577 12552 1582 12608
rect 1638 12552 2084 12608
rect 1577 12550 2084 12552
rect 1577 12547 1643 12550
rect 2078 12548 2084 12550
rect 2148 12548 2154 12612
rect 3233 12610 3299 12613
rect 3877 12610 3943 12613
rect 3233 12608 3943 12610
rect 3233 12552 3238 12608
rect 3294 12552 3882 12608
rect 3938 12552 3943 12608
rect 3233 12550 3943 12552
rect 3233 12547 3299 12550
rect 3877 12547 3943 12550
rect 5717 12610 5783 12613
rect 5942 12610 5948 12612
rect 5717 12608 5948 12610
rect 5717 12552 5722 12608
rect 5778 12552 5948 12608
rect 5717 12550 5948 12552
rect 5717 12547 5783 12550
rect 5942 12548 5948 12550
rect 6012 12548 6018 12612
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 1025 12338 1091 12341
rect 5165 12338 5231 12341
rect 1025 12336 5231 12338
rect 1025 12280 1030 12336
rect 1086 12280 5170 12336
rect 5226 12280 5231 12336
rect 1025 12278 5231 12280
rect 1025 12275 1091 12278
rect 5165 12275 5231 12278
rect 3785 12202 3851 12205
rect 3918 12202 3924 12204
rect 3785 12200 3924 12202
rect 3785 12144 3790 12200
rect 3846 12144 3924 12200
rect 3785 12142 3924 12144
rect 3785 12139 3851 12142
rect 3918 12140 3924 12142
rect 3988 12140 3994 12204
rect 7046 12202 7052 12204
rect 4110 12142 7052 12202
rect 0 12066 800 12096
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 0 11976 800 12006
rect 933 12003 999 12006
rect 3049 12066 3115 12069
rect 4110 12066 4170 12142
rect 7046 12140 7052 12142
rect 7116 12140 7122 12204
rect 14365 12202 14431 12205
rect 14365 12200 15210 12202
rect 14365 12144 14370 12200
rect 14426 12144 15210 12200
rect 14365 12142 15210 12144
rect 14365 12139 14431 12142
rect 3049 12064 4170 12066
rect 3049 12008 3054 12064
rect 3110 12008 4170 12064
rect 3049 12006 4170 12008
rect 15150 12096 15210 12142
rect 15150 12006 16000 12096
rect 3049 12003 3115 12006
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 15200 11976 16000 12006
rect 14653 11935 14969 11936
rect 5257 11794 5323 11797
rect 6913 11794 6979 11797
rect 5257 11792 6979 11794
rect 5257 11736 5262 11792
rect 5318 11736 6918 11792
rect 6974 11736 6979 11792
rect 5257 11734 6979 11736
rect 5257 11731 5323 11734
rect 6913 11731 6979 11734
rect 2037 11658 2103 11661
rect 4245 11658 4311 11661
rect 2037 11656 4311 11658
rect 2037 11600 2042 11656
rect 2098 11600 4250 11656
rect 4306 11600 4311 11656
rect 2037 11598 4311 11600
rect 2037 11595 2103 11598
rect 4245 11595 4311 11598
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 12940 11391 13256 11392
rect 0 11250 800 11280
rect 4061 11250 4127 11253
rect 0 11248 4127 11250
rect 0 11192 4066 11248
rect 4122 11192 4127 11248
rect 0 11190 4127 11192
rect 0 11160 800 11190
rect 4061 11187 4127 11190
rect 7097 11250 7163 11253
rect 12566 11250 12572 11252
rect 7097 11248 12572 11250
rect 7097 11192 7102 11248
rect 7158 11192 12572 11248
rect 7097 11190 12572 11192
rect 7097 11187 7163 11190
rect 12566 11188 12572 11190
rect 12636 11188 12642 11252
rect 14365 11250 14431 11253
rect 15200 11250 16000 11280
rect 14365 11248 16000 11250
rect 14365 11192 14370 11248
rect 14426 11192 16000 11248
rect 14365 11190 16000 11192
rect 14365 11187 14431 11190
rect 15200 11160 16000 11190
rect 1342 11052 1348 11116
rect 1412 11114 1418 11116
rect 1669 11114 1735 11117
rect 1412 11112 1735 11114
rect 1412 11056 1674 11112
rect 1730 11056 1735 11112
rect 1412 11054 1735 11056
rect 1412 11052 1418 11054
rect 1669 11051 1735 11054
rect 3049 11114 3115 11117
rect 8477 11114 8543 11117
rect 3049 11112 8543 11114
rect 3049 11056 3054 11112
rect 3110 11056 8482 11112
rect 8538 11056 8543 11112
rect 3049 11054 8543 11056
rect 3049 11051 3115 11054
rect 8477 11051 8543 11054
rect 11789 11114 11855 11117
rect 12750 11114 12756 11116
rect 11789 11112 12756 11114
rect 11789 11056 11794 11112
rect 11850 11056 12756 11112
rect 11789 11054 12756 11056
rect 11789 11051 11855 11054
rect 12750 11052 12756 11054
rect 12820 11052 12826 11116
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 790 10780 796 10844
rect 860 10842 866 10844
rect 2313 10842 2379 10845
rect 860 10840 2379 10842
rect 860 10784 2318 10840
rect 2374 10784 2379 10840
rect 860 10782 2379 10784
rect 860 10780 866 10782
rect 2313 10779 2379 10782
rect 3785 10842 3851 10845
rect 3785 10840 3986 10842
rect 3785 10784 3790 10840
rect 3846 10784 3986 10840
rect 3785 10782 3986 10784
rect 3785 10779 3851 10782
rect 1853 10706 1919 10709
rect 3926 10706 3986 10782
rect 4061 10706 4127 10709
rect 1853 10704 3618 10706
rect 1853 10648 1858 10704
rect 1914 10648 3618 10704
rect 1853 10646 3618 10648
rect 3926 10704 4127 10706
rect 3926 10648 4066 10704
rect 4122 10648 4127 10704
rect 3926 10646 4127 10648
rect 1853 10643 1919 10646
rect 2313 10570 2379 10573
rect 3558 10570 3618 10646
rect 4061 10643 4127 10646
rect 4838 10644 4844 10708
rect 4908 10644 4914 10708
rect 4846 10570 4906 10644
rect 10174 10570 10180 10572
rect 2313 10568 3434 10570
rect 2313 10512 2318 10568
rect 2374 10512 3434 10568
rect 2313 10510 3434 10512
rect 3558 10510 4906 10570
rect 5030 10510 10180 10570
rect 2313 10507 2379 10510
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 3374 10434 3434 10510
rect 5030 10434 5090 10510
rect 10174 10508 10180 10510
rect 10244 10508 10250 10572
rect 13169 10570 13235 10573
rect 14181 10570 14247 10573
rect 13169 10568 14247 10570
rect 13169 10512 13174 10568
rect 13230 10512 14186 10568
rect 14242 10512 14247 10568
rect 13169 10510 14247 10512
rect 13169 10507 13235 10510
rect 14181 10507 14247 10510
rect 3374 10374 5090 10434
rect 14365 10434 14431 10437
rect 15200 10434 16000 10464
rect 14365 10432 16000 10434
rect 14365 10376 14370 10432
rect 14426 10376 16000 10432
rect 14365 10374 16000 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 14365 10371 14431 10374
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 15200 10344 16000 10374
rect 12940 10303 13256 10304
rect 4889 10298 4955 10301
rect 4889 10296 5320 10298
rect 4889 10240 4894 10296
rect 4950 10240 5320 10296
rect 4889 10238 5320 10240
rect 4889 10235 4955 10238
rect 5260 10162 5320 10238
rect 5390 10236 5396 10300
rect 5460 10298 5466 10300
rect 5625 10298 5691 10301
rect 5460 10296 5691 10298
rect 5460 10240 5630 10296
rect 5686 10240 5691 10296
rect 5460 10238 5691 10240
rect 5460 10236 5466 10238
rect 5625 10235 5691 10238
rect 6545 10162 6611 10165
rect 5260 10160 6611 10162
rect 5260 10104 6550 10160
rect 6606 10104 6611 10160
rect 5260 10102 6611 10104
rect 6545 10099 6611 10102
rect 10041 10162 10107 10165
rect 10358 10162 10364 10164
rect 10041 10160 10364 10162
rect 10041 10104 10046 10160
rect 10102 10104 10364 10160
rect 10041 10102 10364 10104
rect 10041 10099 10107 10102
rect 10358 10100 10364 10102
rect 10428 10100 10434 10164
rect 9029 10026 9095 10029
rect 13169 10026 13235 10029
rect 9029 10024 13235 10026
rect 9029 9968 9034 10024
rect 9090 9968 13174 10024
rect 13230 9968 13235 10024
rect 9029 9966 13235 9968
rect 9029 9963 9095 9966
rect 13169 9963 13235 9966
rect 2262 9828 2268 9892
rect 2332 9890 2338 9892
rect 3417 9890 3483 9893
rect 2332 9888 3483 9890
rect 2332 9832 3422 9888
rect 3478 9832 3483 9888
rect 2332 9830 3483 9832
rect 2332 9828 2338 9830
rect 3417 9827 3483 9830
rect 9949 9890 10015 9893
rect 10593 9890 10659 9893
rect 9949 9888 10659 9890
rect 9949 9832 9954 9888
rect 10010 9832 10598 9888
rect 10654 9832 10659 9888
rect 9949 9830 10659 9832
rect 9949 9827 10015 9830
rect 10593 9827 10659 9830
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 14653 9759 14969 9760
rect 0 9618 800 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 9949 9618 10015 9621
rect 10409 9618 10475 9621
rect 9949 9616 10475 9618
rect 9949 9560 9954 9616
rect 10010 9560 10414 9616
rect 10470 9560 10475 9616
rect 9949 9558 10475 9560
rect 9949 9555 10015 9558
rect 10409 9555 10475 9558
rect 14089 9618 14155 9621
rect 15200 9618 16000 9648
rect 14089 9616 16000 9618
rect 14089 9560 14094 9616
rect 14150 9560 16000 9616
rect 14089 9558 16000 9560
rect 14089 9555 14155 9558
rect 15200 9528 16000 9558
rect 2313 9482 2379 9485
rect 3550 9482 3556 9484
rect 2313 9480 3556 9482
rect 2313 9424 2318 9480
rect 2374 9424 3556 9480
rect 2313 9422 3556 9424
rect 2313 9419 2379 9422
rect 3550 9420 3556 9422
rect 3620 9482 3626 9484
rect 12157 9482 12223 9485
rect 3620 9480 12223 9482
rect 3620 9424 12162 9480
rect 12218 9424 12223 9480
rect 3620 9422 12223 9424
rect 3620 9420 3626 9422
rect 12157 9419 12223 9422
rect 3417 9346 3483 9349
rect 5625 9346 5691 9349
rect 3417 9344 5691 9346
rect 3417 9288 3422 9344
rect 3478 9288 5630 9344
rect 5686 9288 5691 9344
rect 3417 9286 5691 9288
rect 3417 9283 3483 9286
rect 5625 9283 5691 9286
rect 10358 9284 10364 9348
rect 10428 9284 10434 9348
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 10366 9210 10426 9284
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 10501 9210 10567 9213
rect 10366 9208 10567 9210
rect 10366 9152 10506 9208
rect 10562 9152 10567 9208
rect 10366 9150 10567 9152
rect 10501 9147 10567 9150
rect 2221 9074 2287 9077
rect 3182 9074 3188 9076
rect 2221 9072 3188 9074
rect 2221 9016 2226 9072
rect 2282 9016 3188 9072
rect 2221 9014 3188 9016
rect 2221 9011 2287 9014
rect 3182 9012 3188 9014
rect 3252 9012 3258 9076
rect 4705 9074 4771 9077
rect 6862 9074 6868 9076
rect 4705 9072 6868 9074
rect 4705 9016 4710 9072
rect 4766 9016 6868 9072
rect 4705 9014 6868 9016
rect 4705 9011 4771 9014
rect 6862 9012 6868 9014
rect 6932 9012 6938 9076
rect 3734 8876 3740 8940
rect 3804 8938 3810 8940
rect 7925 8938 7991 8941
rect 3804 8936 7991 8938
rect 3804 8880 7930 8936
rect 7986 8880 7991 8936
rect 3804 8878 7991 8880
rect 3804 8876 3810 8878
rect 7925 8875 7991 8878
rect 14365 8938 14431 8941
rect 14365 8936 15210 8938
rect 14365 8880 14370 8936
rect 14426 8880 15210 8936
rect 14365 8878 15210 8880
rect 14365 8875 14431 8878
rect 15150 8832 15210 8878
rect 0 8802 800 8832
rect 0 8742 1042 8802
rect 15150 8742 16000 8832
rect 0 8712 800 8742
rect 982 8394 1042 8742
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 15200 8712 16000 8742
rect 14653 8671 14969 8672
rect 11697 8666 11763 8669
rect 13537 8666 13603 8669
rect 11697 8664 13603 8666
rect 11697 8608 11702 8664
rect 11758 8608 13542 8664
rect 13598 8608 13603 8664
rect 11697 8606 13603 8608
rect 11697 8603 11763 8606
rect 13537 8603 13603 8606
rect 4705 8530 4771 8533
rect 9489 8530 9555 8533
rect 3742 8528 4771 8530
rect 3742 8472 4710 8528
rect 4766 8472 4771 8528
rect 3742 8470 4771 8472
rect 1853 8394 1919 8397
rect 982 8392 1919 8394
rect 982 8336 1858 8392
rect 1914 8336 1919 8392
rect 982 8334 1919 8336
rect 1853 8331 1919 8334
rect 2446 8332 2452 8396
rect 2516 8394 2522 8396
rect 2589 8394 2655 8397
rect 2516 8392 2655 8394
rect 2516 8336 2594 8392
rect 2650 8336 2655 8392
rect 2516 8334 2655 8336
rect 2516 8332 2522 8334
rect 2589 8331 2655 8334
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 0 7986 800 8016
rect 1485 7986 1551 7989
rect 1894 7986 1900 7988
rect 0 7926 1410 7986
rect 0 7896 800 7926
rect 1350 7714 1410 7926
rect 1485 7984 1900 7986
rect 1485 7928 1490 7984
rect 1546 7928 1900 7984
rect 1485 7926 1900 7928
rect 1485 7923 1551 7926
rect 1894 7924 1900 7926
rect 1964 7924 1970 7988
rect 2313 7986 2379 7989
rect 3742 7986 3802 8470
rect 4705 8467 4771 8470
rect 9262 8528 9555 8530
rect 9262 8472 9494 8528
rect 9550 8472 9555 8528
rect 9262 8470 9555 8472
rect 8518 8196 8524 8260
rect 8588 8258 8594 8260
rect 8845 8258 8911 8261
rect 8588 8256 8911 8258
rect 8588 8200 8850 8256
rect 8906 8200 8911 8256
rect 8588 8198 8911 8200
rect 8588 8196 8594 8198
rect 8845 8195 8911 8198
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 4429 8122 4495 8125
rect 5901 8122 5967 8125
rect 4429 8120 5967 8122
rect 4429 8064 4434 8120
rect 4490 8064 5906 8120
rect 5962 8064 5967 8120
rect 4429 8062 5967 8064
rect 4429 8059 4495 8062
rect 5901 8059 5967 8062
rect 9262 7989 9322 8470
rect 9489 8467 9555 8470
rect 10358 8468 10364 8532
rect 10428 8530 10434 8532
rect 10869 8530 10935 8533
rect 10428 8528 10935 8530
rect 10428 8472 10874 8528
rect 10930 8472 10935 8528
rect 10428 8470 10935 8472
rect 10428 8468 10434 8470
rect 10869 8467 10935 8470
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 12940 8127 13256 8128
rect 2313 7984 3802 7986
rect 2313 7928 2318 7984
rect 2374 7928 3802 7984
rect 2313 7926 3802 7928
rect 5441 7986 5507 7989
rect 6678 7986 6684 7988
rect 5441 7984 6684 7986
rect 5441 7928 5446 7984
rect 5502 7928 6684 7984
rect 5441 7926 6684 7928
rect 2313 7923 2379 7926
rect 5441 7923 5507 7926
rect 6678 7924 6684 7926
rect 6748 7924 6754 7988
rect 9262 7984 9371 7989
rect 9262 7928 9310 7984
rect 9366 7928 9371 7984
rect 9262 7926 9371 7928
rect 9305 7923 9371 7926
rect 11697 7986 11763 7989
rect 15200 7986 16000 8016
rect 11697 7984 16000 7986
rect 11697 7928 11702 7984
rect 11758 7928 16000 7984
rect 11697 7926 16000 7928
rect 11697 7923 11763 7926
rect 15200 7896 16000 7926
rect 1485 7850 1551 7853
rect 8569 7850 8635 7853
rect 1485 7848 8635 7850
rect 1485 7792 1490 7848
rect 1546 7792 8574 7848
rect 8630 7792 8635 7848
rect 1485 7790 8635 7792
rect 1485 7787 1551 7790
rect 8569 7787 8635 7790
rect 10726 7788 10732 7852
rect 10796 7850 10802 7852
rect 11329 7850 11395 7853
rect 10796 7848 11395 7850
rect 10796 7792 11334 7848
rect 11390 7792 11395 7848
rect 10796 7790 11395 7792
rect 10796 7788 10802 7790
rect 11329 7787 11395 7790
rect 3969 7714 4035 7717
rect 1350 7712 4035 7714
rect 1350 7656 3974 7712
rect 4030 7656 4035 7712
rect 1350 7654 4035 7656
rect 3969 7651 4035 7654
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 5073 7442 5139 7445
rect 1350 7440 5139 7442
rect 1350 7384 5078 7440
rect 5134 7384 5139 7440
rect 1350 7382 5139 7384
rect 0 7170 800 7200
rect 1350 7170 1410 7382
rect 5073 7379 5139 7382
rect 1485 7306 1551 7309
rect 10961 7308 11027 7309
rect 2262 7306 2268 7308
rect 1485 7304 2268 7306
rect 1485 7248 1490 7304
rect 1546 7248 2268 7304
rect 1485 7246 2268 7248
rect 1485 7243 1551 7246
rect 2262 7244 2268 7246
rect 2332 7244 2338 7308
rect 10910 7306 10916 7308
rect 10870 7246 10916 7306
rect 10980 7304 11027 7308
rect 11022 7248 11027 7304
rect 10910 7244 10916 7246
rect 10980 7244 11027 7248
rect 10961 7243 11027 7244
rect 0 7110 1410 7170
rect 13721 7170 13787 7173
rect 15200 7170 16000 7200
rect 13721 7168 16000 7170
rect 13721 7112 13726 7168
rect 13782 7112 16000 7168
rect 13721 7110 16000 7112
rect 0 7080 800 7110
rect 13721 7107 13787 7110
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 15200 7080 16000 7110
rect 12940 7039 13256 7040
rect 3877 7036 3943 7037
rect 3877 7034 3924 7036
rect 3832 7032 3924 7034
rect 3832 6976 3882 7032
rect 3832 6974 3924 6976
rect 3877 6972 3924 6974
rect 3988 6972 3994 7036
rect 3877 6971 3943 6972
rect 2037 6900 2103 6901
rect 2037 6896 2084 6900
rect 2148 6898 2154 6900
rect 2037 6840 2042 6896
rect 2037 6836 2084 6840
rect 2148 6838 2194 6898
rect 2148 6836 2154 6838
rect 2037 6835 2103 6836
rect 11145 6762 11211 6765
rect 11145 6760 11714 6762
rect 11145 6704 11150 6760
rect 11206 6704 11714 6760
rect 11145 6702 11714 6704
rect 11145 6699 11211 6702
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 0 6354 800 6384
rect 11654 6357 11714 6702
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 12617 6492 12683 6493
rect 12566 6428 12572 6492
rect 12636 6490 12683 6492
rect 12636 6488 12728 6490
rect 12678 6432 12728 6488
rect 12636 6430 12728 6432
rect 12636 6428 12683 6430
rect 12617 6427 12683 6428
rect 1393 6354 1459 6357
rect 0 6352 1459 6354
rect 0 6296 1398 6352
rect 1454 6296 1459 6352
rect 0 6294 1459 6296
rect 0 6264 800 6294
rect 1393 6291 1459 6294
rect 4613 6354 4679 6357
rect 8334 6354 8340 6356
rect 4613 6352 8340 6354
rect 4613 6296 4618 6352
rect 4674 6296 8340 6352
rect 4613 6294 8340 6296
rect 4613 6291 4679 6294
rect 8334 6292 8340 6294
rect 8404 6292 8410 6356
rect 11654 6352 11763 6357
rect 11654 6296 11702 6352
rect 11758 6296 11763 6352
rect 11654 6294 11763 6296
rect 11697 6291 11763 6294
rect 12249 6354 12315 6357
rect 15200 6354 16000 6384
rect 12249 6352 16000 6354
rect 12249 6296 12254 6352
rect 12310 6296 16000 6352
rect 12249 6294 16000 6296
rect 12249 6291 12315 6294
rect 15200 6264 16000 6294
rect 3366 6156 3372 6220
rect 3436 6218 3442 6220
rect 9489 6218 9555 6221
rect 3436 6216 9555 6218
rect 3436 6160 9494 6216
rect 9550 6160 9555 6216
rect 3436 6158 9555 6160
rect 3436 6156 3442 6158
rect 9489 6155 9555 6158
rect 3969 6082 4035 6085
rect 5165 6082 5231 6085
rect 3969 6080 5231 6082
rect 3969 6024 3974 6080
rect 4030 6024 5170 6080
rect 5226 6024 5231 6080
rect 3969 6022 5231 6024
rect 3969 6019 4035 6022
rect 5165 6019 5231 6022
rect 7097 6082 7163 6085
rect 8845 6082 8911 6085
rect 7097 6080 8911 6082
rect 7097 6024 7102 6080
rect 7158 6024 8850 6080
rect 8906 6024 8911 6080
rect 7097 6022 8911 6024
rect 7097 6019 7163 6022
rect 8845 6019 8911 6022
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 6361 5810 6427 5813
rect 11237 5810 11303 5813
rect 6361 5808 11303 5810
rect 6361 5752 6366 5808
rect 6422 5752 11242 5808
rect 11298 5752 11303 5808
rect 6361 5750 11303 5752
rect 6361 5747 6427 5750
rect 11237 5747 11303 5750
rect 5809 5674 5875 5677
rect 8201 5674 8267 5677
rect 5809 5672 8267 5674
rect 5809 5616 5814 5672
rect 5870 5616 8206 5672
rect 8262 5616 8267 5672
rect 5809 5614 8267 5616
rect 5809 5611 5875 5614
rect 8201 5611 8267 5614
rect 10777 5674 10843 5677
rect 12341 5674 12407 5677
rect 10777 5672 12407 5674
rect 10777 5616 10782 5672
rect 10838 5616 12346 5672
rect 12402 5616 12407 5672
rect 10777 5614 12407 5616
rect 10777 5611 10843 5614
rect 12341 5611 12407 5614
rect 0 5538 800 5568
rect 1669 5538 1735 5541
rect 15200 5538 16000 5568
rect 0 5536 1735 5538
rect 0 5480 1674 5536
rect 1730 5480 1735 5536
rect 0 5478 1735 5480
rect 0 5448 800 5478
rect 1669 5475 1735 5478
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 15150 5448 16000 5538
rect 6177 5402 6243 5405
rect 11973 5402 12039 5405
rect 4892 5400 6243 5402
rect 4892 5344 6182 5400
rect 6238 5344 6243 5400
rect 4892 5342 6243 5344
rect 1301 5266 1367 5269
rect 4892 5266 4952 5342
rect 6177 5339 6243 5342
rect 11654 5400 12039 5402
rect 11654 5344 11978 5400
rect 12034 5344 12039 5400
rect 11654 5342 12039 5344
rect 1301 5264 4952 5266
rect 1301 5208 1306 5264
rect 1362 5208 4952 5264
rect 1301 5206 4952 5208
rect 5073 5266 5139 5269
rect 11654 5266 11714 5342
rect 11973 5339 12039 5342
rect 5073 5264 11714 5266
rect 5073 5208 5078 5264
rect 5134 5208 11714 5264
rect 5073 5206 11714 5208
rect 1301 5203 1367 5206
rect 5073 5203 5139 5206
rect 3509 5130 3575 5133
rect 6085 5130 6151 5133
rect 3509 5128 6151 5130
rect 3509 5072 3514 5128
rect 3570 5072 6090 5128
rect 6146 5072 6151 5128
rect 3509 5070 6151 5072
rect 3509 5067 3575 5070
rect 6085 5067 6151 5070
rect 6821 5130 6887 5133
rect 8569 5130 8635 5133
rect 10685 5130 10751 5133
rect 15150 5130 15210 5448
rect 6821 5128 8635 5130
rect 6821 5072 6826 5128
rect 6882 5072 8574 5128
rect 8630 5072 8635 5128
rect 6821 5070 8635 5072
rect 6821 5067 6887 5070
rect 8569 5067 8635 5070
rect 9262 5128 10751 5130
rect 9262 5072 10690 5128
rect 10746 5072 10751 5128
rect 9262 5070 10751 5072
rect 6545 4994 6611 4997
rect 9262 4994 9322 5070
rect 10685 5067 10751 5070
rect 12390 5070 15210 5130
rect 6545 4992 9322 4994
rect 6545 4936 6550 4992
rect 6606 4936 9322 4992
rect 6545 4934 9322 4936
rect 6545 4931 6611 4934
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 6678 4796 6684 4860
rect 6748 4858 6754 4860
rect 6913 4858 6979 4861
rect 6748 4856 6979 4858
rect 6748 4800 6918 4856
rect 6974 4800 6979 4856
rect 6748 4798 6979 4800
rect 6748 4796 6754 4798
rect 6913 4795 6979 4798
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 5349 4722 5415 4725
rect 9990 4722 9996 4724
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 3190 4720 5415 4722
rect 3190 4664 5354 4720
rect 5410 4664 5415 4720
rect 3190 4662 5415 4664
rect 1945 4586 2011 4589
rect 3190 4586 3250 4662
rect 5349 4659 5415 4662
rect 9630 4662 9996 4722
rect 1945 4584 3250 4586
rect 1945 4528 1950 4584
rect 2006 4528 3250 4584
rect 1945 4526 3250 4528
rect 1945 4523 2011 4526
rect 3918 4524 3924 4588
rect 3988 4586 3994 4588
rect 9630 4586 9690 4662
rect 9990 4660 9996 4662
rect 10060 4722 10066 4724
rect 12390 4722 12450 5070
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 12940 4863 13256 4864
rect 10060 4662 12450 4722
rect 13721 4722 13787 4725
rect 15200 4722 16000 4752
rect 13721 4720 16000 4722
rect 13721 4664 13726 4720
rect 13782 4664 16000 4720
rect 13721 4662 16000 4664
rect 10060 4660 10066 4662
rect 13721 4659 13787 4662
rect 15200 4632 16000 4662
rect 3988 4526 9690 4586
rect 9857 4586 9923 4589
rect 10685 4586 10751 4589
rect 13445 4586 13511 4589
rect 9857 4584 13511 4586
rect 9857 4528 9862 4584
rect 9918 4528 10690 4584
rect 10746 4528 13450 4584
rect 13506 4528 13511 4584
rect 9857 4526 13511 4528
rect 3988 4524 3994 4526
rect 9857 4523 9923 4526
rect 10685 4523 10751 4526
rect 13445 4523 13511 4526
rect 4889 4450 4955 4453
rect 6545 4450 6611 4453
rect 4889 4448 6611 4450
rect 4889 4392 4894 4448
rect 4950 4392 6550 4448
rect 6606 4392 6611 4448
rect 4889 4390 6611 4392
rect 4889 4387 4955 4390
rect 6545 4387 6611 4390
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 5717 4314 5783 4317
rect 6361 4314 6427 4317
rect 5717 4312 6427 4314
rect 5717 4256 5722 4312
rect 5778 4256 6366 4312
rect 6422 4256 6427 4312
rect 5717 4254 6427 4256
rect 5717 4251 5783 4254
rect 6361 4251 6427 4254
rect 9990 4252 9996 4316
rect 10060 4314 10066 4316
rect 10317 4314 10383 4317
rect 10060 4312 10383 4314
rect 10060 4256 10322 4312
rect 10378 4256 10383 4312
rect 10060 4254 10383 4256
rect 10060 4252 10066 4254
rect 10317 4251 10383 4254
rect 2221 4178 2287 4181
rect 3734 4178 3740 4180
rect 2221 4176 3740 4178
rect 2221 4120 2226 4176
rect 2282 4120 3740 4176
rect 2221 4118 3740 4120
rect 2221 4115 2287 4118
rect 3734 4116 3740 4118
rect 3804 4116 3810 4180
rect 4061 4178 4127 4181
rect 11973 4178 12039 4181
rect 4061 4176 12039 4178
rect 4061 4120 4066 4176
rect 4122 4120 11978 4176
rect 12034 4120 12039 4176
rect 4061 4118 12039 4120
rect 4061 4115 4127 4118
rect 11973 4115 12039 4118
rect 1894 3980 1900 4044
rect 1964 4042 1970 4044
rect 2405 4042 2471 4045
rect 1964 4040 2471 4042
rect 1964 3984 2410 4040
rect 2466 3984 2471 4040
rect 1964 3982 2471 3984
rect 1964 3980 1970 3982
rect 2405 3979 2471 3982
rect 2957 4042 3023 4045
rect 4797 4042 4863 4045
rect 5390 4042 5396 4044
rect 2957 4040 5396 4042
rect 2957 3984 2962 4040
rect 3018 3984 4802 4040
rect 4858 3984 5396 4040
rect 2957 3982 5396 3984
rect 2957 3979 3023 3982
rect 4797 3979 4863 3982
rect 5390 3980 5396 3982
rect 5460 3980 5466 4044
rect 5574 3980 5580 4044
rect 5644 4042 5650 4044
rect 5993 4042 6059 4045
rect 5644 4040 6059 4042
rect 5644 3984 5998 4040
rect 6054 3984 6059 4040
rect 5644 3982 6059 3984
rect 5644 3980 5650 3982
rect 5993 3979 6059 3982
rect 6494 3980 6500 4044
rect 6564 4042 6570 4044
rect 8385 4042 8451 4045
rect 6564 4040 8451 4042
rect 6564 3984 8390 4040
rect 8446 3984 8451 4040
rect 6564 3982 8451 3984
rect 6564 3980 6570 3982
rect 8385 3979 8451 3982
rect 10910 3980 10916 4044
rect 10980 3980 10986 4044
rect 0 3906 800 3936
rect 3325 3906 3391 3909
rect 5257 3906 5323 3909
rect 0 3846 1410 3906
rect 0 3816 800 3846
rect 1350 3634 1410 3846
rect 3325 3904 5323 3906
rect 3325 3848 3330 3904
rect 3386 3848 5262 3904
rect 5318 3848 5323 3904
rect 3325 3846 5323 3848
rect 3325 3843 3391 3846
rect 5257 3843 5323 3846
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 3785 3770 3851 3773
rect 5717 3770 5783 3773
rect 5942 3770 5948 3772
rect 3785 3768 5948 3770
rect 3785 3712 3790 3768
rect 3846 3712 5722 3768
rect 5778 3712 5948 3768
rect 3785 3710 5948 3712
rect 3785 3707 3851 3710
rect 5717 3707 5783 3710
rect 5942 3708 5948 3710
rect 6012 3708 6018 3772
rect 3877 3634 3943 3637
rect 1350 3632 3943 3634
rect 1350 3576 3882 3632
rect 3938 3576 3943 3632
rect 1350 3574 3943 3576
rect 3877 3571 3943 3574
rect 5625 3634 5691 3637
rect 10918 3634 10978 3980
rect 15200 3906 16000 3936
rect 13448 3846 16000 3906
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 11053 3770 11119 3773
rect 11053 3768 11530 3770
rect 11053 3712 11058 3768
rect 11114 3712 11530 3768
rect 11053 3710 11530 3712
rect 11053 3707 11119 3710
rect 5625 3632 10978 3634
rect 5625 3576 5630 3632
rect 5686 3576 10978 3632
rect 5625 3574 10978 3576
rect 11470 3634 11530 3710
rect 11605 3634 11671 3637
rect 11470 3632 11671 3634
rect 11470 3576 11610 3632
rect 11666 3576 11671 3632
rect 11470 3574 11671 3576
rect 5625 3571 5691 3574
rect 11605 3571 11671 3574
rect 12157 3634 12223 3637
rect 13448 3634 13508 3846
rect 15200 3816 16000 3846
rect 12157 3632 13508 3634
rect 12157 3576 12162 3632
rect 12218 3576 13508 3632
rect 12157 3574 13508 3576
rect 12157 3571 12223 3574
rect 974 3436 980 3500
rect 1044 3498 1050 3500
rect 3233 3498 3299 3501
rect 1044 3496 3299 3498
rect 1044 3440 3238 3496
rect 3294 3440 3299 3496
rect 1044 3438 3299 3440
rect 1044 3436 1050 3438
rect 3233 3435 3299 3438
rect 3550 3436 3556 3500
rect 3620 3498 3626 3500
rect 3877 3498 3943 3501
rect 6545 3498 6611 3501
rect 11329 3498 11395 3501
rect 3620 3496 3943 3498
rect 3620 3440 3882 3496
rect 3938 3440 3943 3496
rect 3620 3438 3943 3440
rect 3620 3436 3626 3438
rect 3877 3435 3943 3438
rect 4248 3496 6611 3498
rect 4248 3440 6550 3496
rect 6606 3440 6611 3496
rect 4248 3438 6611 3440
rect 565 3362 631 3365
rect 3233 3364 3299 3365
rect 565 3360 2790 3362
rect 565 3304 570 3360
rect 626 3304 2790 3360
rect 565 3302 2790 3304
rect 565 3299 631 3302
rect 0 3090 800 3120
rect 1342 3090 1348 3092
rect 0 3030 1348 3090
rect 0 3000 800 3030
rect 1342 3028 1348 3030
rect 1412 3028 1418 3092
rect 2730 3090 2790 3302
rect 3182 3300 3188 3364
rect 3252 3362 3299 3364
rect 4248 3362 4308 3438
rect 6545 3435 6611 3438
rect 6686 3496 11395 3498
rect 6686 3440 11334 3496
rect 11390 3440 11395 3496
rect 6686 3438 11395 3440
rect 3252 3360 4308 3362
rect 3294 3304 4308 3360
rect 3252 3302 4308 3304
rect 5717 3362 5783 3365
rect 6686 3362 6746 3438
rect 11329 3435 11395 3438
rect 5717 3360 6746 3362
rect 5717 3304 5722 3360
rect 5778 3304 6746 3360
rect 5717 3302 6746 3304
rect 8385 3362 8451 3365
rect 10869 3362 10935 3365
rect 12341 3362 12407 3365
rect 8385 3360 10935 3362
rect 8385 3304 8390 3360
rect 8446 3304 10874 3360
rect 10930 3304 10935 3360
rect 8385 3302 10935 3304
rect 3252 3300 3299 3302
rect 3233 3299 3299 3300
rect 5717 3299 5783 3302
rect 8385 3299 8451 3302
rect 10869 3299 10935 3302
rect 11654 3360 12407 3362
rect 11654 3304 12346 3360
rect 12402 3304 12407 3360
rect 11654 3302 12407 3304
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 6862 3164 6868 3228
rect 6932 3226 6938 3228
rect 7649 3226 7715 3229
rect 6932 3224 7715 3226
rect 6932 3168 7654 3224
rect 7710 3168 7715 3224
rect 6932 3166 7715 3168
rect 6932 3164 6938 3166
rect 7649 3163 7715 3166
rect 4981 3090 5047 3093
rect 2730 3088 5047 3090
rect 2730 3032 4986 3088
rect 5042 3032 5047 3088
rect 2730 3030 5047 3032
rect 4981 3027 5047 3030
rect 7414 3028 7420 3092
rect 7484 3090 7490 3092
rect 7925 3090 7991 3093
rect 7484 3088 7991 3090
rect 7484 3032 7930 3088
rect 7986 3032 7991 3088
rect 7484 3030 7991 3032
rect 7484 3028 7490 3030
rect 7925 3027 7991 3030
rect 1485 2954 1551 2957
rect 11654 2954 11714 3302
rect 12341 3299 12407 3302
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 14457 3090 14523 3093
rect 15200 3090 16000 3120
rect 14457 3088 16000 3090
rect 14457 3032 14462 3088
rect 14518 3032 16000 3088
rect 14457 3030 16000 3032
rect 14457 3027 14523 3030
rect 15200 3000 16000 3030
rect 1485 2952 11714 2954
rect 1485 2896 1490 2952
rect 1546 2896 11714 2952
rect 1485 2894 11714 2896
rect 12525 2954 12591 2957
rect 12750 2954 12756 2956
rect 12525 2952 12756 2954
rect 12525 2896 12530 2952
rect 12586 2896 12756 2952
rect 12525 2894 12756 2896
rect 1485 2891 1551 2894
rect 12525 2891 12591 2894
rect 12750 2892 12756 2894
rect 12820 2892 12826 2956
rect 4245 2818 4311 2821
rect 4838 2818 4844 2820
rect 4245 2816 4844 2818
rect 4245 2760 4250 2816
rect 4306 2760 4844 2816
rect 4245 2758 4844 2760
rect 4245 2755 4311 2758
rect 4838 2756 4844 2758
rect 4908 2756 4914 2820
rect 6494 2756 6500 2820
rect 6564 2756 6570 2820
rect 7046 2756 7052 2820
rect 7116 2818 7122 2820
rect 7741 2818 7807 2821
rect 7116 2816 7807 2818
rect 7116 2760 7746 2816
rect 7802 2760 7807 2816
rect 7116 2758 7807 2760
rect 7116 2756 7122 2758
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 3141 2682 3207 2685
rect 3366 2682 3372 2684
rect 3141 2680 3372 2682
rect 3141 2624 3146 2680
rect 3202 2624 3372 2680
rect 3141 2622 3372 2624
rect 3141 2619 3207 2622
rect 3366 2620 3372 2622
rect 3436 2620 3442 2684
rect 4102 2620 4108 2684
rect 4172 2682 4178 2684
rect 4613 2682 4679 2685
rect 4172 2680 4679 2682
rect 4172 2624 4618 2680
rect 4674 2624 4679 2680
rect 4172 2622 4679 2624
rect 4172 2620 4178 2622
rect 4613 2619 4679 2622
rect 2589 2546 2655 2549
rect 3918 2546 3924 2548
rect 2589 2544 3924 2546
rect 2589 2488 2594 2544
rect 2650 2488 3924 2544
rect 2589 2486 3924 2488
rect 2589 2483 2655 2486
rect 3918 2484 3924 2486
rect 3988 2484 3994 2548
rect 4061 2546 4127 2549
rect 6502 2546 6562 2756
rect 7741 2755 7807 2758
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 6637 2682 6703 2685
rect 9213 2682 9279 2685
rect 10777 2684 10843 2685
rect 6637 2680 9279 2682
rect 6637 2624 6642 2680
rect 6698 2624 9218 2680
rect 9274 2624 9279 2680
rect 6637 2622 9279 2624
rect 6637 2619 6703 2622
rect 9213 2619 9279 2622
rect 10358 2620 10364 2684
rect 10428 2620 10434 2684
rect 10726 2620 10732 2684
rect 10796 2682 10843 2684
rect 10796 2680 10888 2682
rect 10838 2624 10888 2680
rect 10796 2622 10888 2624
rect 10796 2620 10843 2622
rect 4061 2544 6562 2546
rect 4061 2488 4066 2544
rect 4122 2488 6562 2544
rect 4061 2486 6562 2488
rect 9029 2548 9095 2549
rect 9029 2544 9076 2548
rect 9140 2546 9146 2548
rect 9765 2546 9831 2549
rect 10225 2546 10291 2549
rect 9029 2488 9034 2544
rect 4061 2483 4127 2486
rect 9029 2484 9076 2488
rect 9140 2486 9186 2546
rect 9765 2544 10291 2546
rect 9765 2488 9770 2544
rect 9826 2488 10230 2544
rect 10286 2488 10291 2544
rect 9765 2486 10291 2488
rect 9140 2484 9146 2486
rect 9029 2483 9095 2484
rect 9765 2483 9831 2486
rect 10225 2483 10291 2486
rect 3325 2410 3391 2413
rect 10366 2410 10426 2620
rect 10777 2619 10843 2620
rect 11881 2546 11947 2549
rect 14273 2546 14339 2549
rect 11881 2544 14339 2546
rect 11881 2488 11886 2544
rect 11942 2488 14278 2544
rect 14334 2488 14339 2544
rect 11881 2486 14339 2488
rect 11881 2483 11947 2486
rect 14273 2483 14339 2486
rect 3325 2408 10426 2410
rect 3325 2352 3330 2408
rect 3386 2352 10426 2408
rect 3325 2350 10426 2352
rect 12065 2410 12131 2413
rect 12065 2408 15210 2410
rect 12065 2352 12070 2408
rect 12126 2352 15210 2408
rect 12065 2350 15210 2352
rect 3325 2347 3391 2350
rect 12065 2347 12131 2350
rect 15150 2304 15210 2350
rect 0 2274 800 2304
rect 0 2214 2790 2274
rect 0 2184 800 2214
rect 2730 2002 2790 2214
rect 10174 2212 10180 2276
rect 10244 2212 10250 2276
rect 15150 2214 16000 2304
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 10182 2002 10242 2212
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 15200 2184 16000 2214
rect 14653 2143 14969 2144
rect 2730 1942 10242 2002
rect 790 1804 796 1868
rect 860 1866 866 1868
rect 5349 1866 5415 1869
rect 860 1864 5415 1866
rect 860 1808 5354 1864
rect 5410 1808 5415 1864
rect 860 1806 5415 1808
rect 860 1804 866 1806
rect 5349 1803 5415 1806
rect 1158 1532 1164 1596
rect 1228 1594 1234 1596
rect 7097 1594 7163 1597
rect 1228 1592 7163 1594
rect 1228 1536 7102 1592
rect 7158 1536 7163 1592
rect 1228 1534 7163 1536
rect 1228 1532 1234 1534
rect 7097 1531 7163 1534
rect 9949 1460 10015 1461
rect 9949 1458 9996 1460
rect 9904 1456 9996 1458
rect 9904 1400 9954 1456
rect 9904 1398 9996 1400
rect 9949 1396 9996 1398
rect 10060 1396 10066 1460
rect 11237 1458 11303 1461
rect 15200 1458 16000 1488
rect 11237 1456 16000 1458
rect 11237 1400 11242 1456
rect 11298 1400 16000 1456
rect 11237 1398 16000 1400
rect 9949 1395 10015 1396
rect 11237 1395 11303 1398
rect 15200 1368 16000 1398
rect 2446 716 2452 780
rect 2516 778 2522 780
rect 2681 778 2747 781
rect 2516 776 2747 778
rect 2516 720 2686 776
rect 2742 720 2747 776
rect 2516 718 2747 720
rect 2516 716 2522 718
rect 2681 715 2747 718
<< via3 >>
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 8340 14452 8404 14516
rect 8524 14316 8588 14380
rect 1164 14180 1228 14244
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 980 13772 1044 13836
rect 9076 13908 9140 13972
rect 9996 13772 10060 13836
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 6500 13092 6564 13156
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 4108 12956 4172 13020
rect 5580 12956 5644 13020
rect 7420 12820 7484 12884
rect 2084 12548 2148 12612
rect 5948 12548 6012 12612
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 3924 12140 3988 12204
rect 7052 12140 7116 12204
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 12572 11188 12636 11252
rect 1348 11052 1412 11116
rect 12756 11052 12820 11116
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 796 10780 860 10844
rect 4844 10644 4908 10708
rect 10180 10508 10244 10572
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 5396 10236 5460 10300
rect 10364 10100 10428 10164
rect 2268 9828 2332 9892
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 3556 9420 3620 9484
rect 10364 9284 10428 9348
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 3188 9012 3252 9076
rect 6868 9012 6932 9076
rect 3740 8876 3804 8940
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2452 8332 2516 8396
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 1900 7924 1964 7988
rect 8524 8196 8588 8260
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 10364 8468 10428 8532
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 6684 7924 6748 7988
rect 10732 7788 10796 7852
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2268 7244 2332 7308
rect 10916 7304 10980 7308
rect 10916 7248 10966 7304
rect 10966 7248 10980 7304
rect 10916 7244 10980 7248
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 3924 7032 3988 7036
rect 3924 6976 3938 7032
rect 3938 6976 3988 7032
rect 3924 6972 3988 6976
rect 2084 6896 2148 6900
rect 2084 6840 2098 6896
rect 2098 6840 2148 6896
rect 2084 6836 2148 6840
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 12572 6488 12636 6492
rect 12572 6432 12622 6488
rect 12622 6432 12636 6488
rect 12572 6428 12636 6432
rect 8340 6292 8404 6356
rect 3372 6156 3436 6220
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 6684 4796 6748 4860
rect 3924 4524 3988 4588
rect 9996 4660 10060 4724
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 9996 4252 10060 4316
rect 3740 4116 3804 4180
rect 1900 3980 1964 4044
rect 5396 3980 5460 4044
rect 5580 3980 5644 4044
rect 6500 3980 6564 4044
rect 10916 3980 10980 4044
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 5948 3708 6012 3772
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 980 3436 1044 3500
rect 3556 3436 3620 3500
rect 1348 3028 1412 3092
rect 3188 3360 3252 3364
rect 3188 3304 3238 3360
rect 3238 3304 3252 3360
rect 3188 3300 3252 3304
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 6868 3164 6932 3228
rect 7420 3028 7484 3092
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 12756 2892 12820 2956
rect 4844 2756 4908 2820
rect 6500 2756 6564 2820
rect 7052 2756 7116 2820
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 3372 2620 3436 2684
rect 4108 2620 4172 2684
rect 3924 2484 3988 2548
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 10364 2620 10428 2684
rect 10732 2680 10796 2684
rect 10732 2624 10782 2680
rect 10782 2624 10796 2680
rect 10732 2620 10796 2624
rect 9076 2544 9140 2548
rect 9076 2488 9090 2544
rect 9090 2488 9140 2544
rect 9076 2484 9140 2488
rect 10180 2212 10244 2276
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
rect 796 1804 860 1868
rect 1164 1532 1228 1596
rect 9996 1456 10060 1460
rect 9996 1400 10010 1456
rect 10010 1400 10060 1456
rect 9996 1396 10060 1400
rect 2452 716 2516 780
<< metal4 >>
rect 2657 16896 2977 17456
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 1163 14244 1229 14245
rect 1163 14180 1164 14244
rect 1228 14180 1229 14244
rect 1163 14179 1229 14180
rect 979 13836 1045 13837
rect 979 13772 980 13836
rect 1044 13772 1045 13836
rect 979 13771 1045 13772
rect 795 10844 861 10845
rect 795 10780 796 10844
rect 860 10780 861 10844
rect 795 10779 861 10780
rect 798 1869 858 10779
rect 982 3501 1042 13771
rect 979 3500 1045 3501
rect 979 3436 980 3500
rect 1044 3436 1045 3500
rect 979 3435 1045 3436
rect 795 1868 861 1869
rect 795 1804 796 1868
rect 860 1804 861 1868
rect 795 1803 861 1804
rect 1166 1597 1226 14179
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2083 12612 2149 12613
rect 2083 12548 2084 12612
rect 2148 12548 2149 12612
rect 2083 12547 2149 12548
rect 1347 11116 1413 11117
rect 1347 11052 1348 11116
rect 1412 11052 1413 11116
rect 1347 11051 1413 11052
rect 1350 3093 1410 11051
rect 1899 7988 1965 7989
rect 1899 7924 1900 7988
rect 1964 7924 1965 7988
rect 1899 7923 1965 7924
rect 1902 4045 1962 7923
rect 2086 6901 2146 12547
rect 2657 12544 2977 13568
rect 4370 17440 4690 17456
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4107 13020 4173 13021
rect 4107 12956 4108 13020
rect 4172 12956 4173 13020
rect 4107 12955 4173 12956
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 3923 12204 3989 12205
rect 3923 12140 3924 12204
rect 3988 12140 3989 12204
rect 3923 12139 3989 12140
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2267 9892 2333 9893
rect 2267 9828 2268 9892
rect 2332 9828 2333 9892
rect 2267 9827 2333 9828
rect 2270 7309 2330 9827
rect 2657 9280 2977 10304
rect 3555 9484 3621 9485
rect 3555 9420 3556 9484
rect 3620 9420 3621 9484
rect 3555 9419 3621 9420
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2451 8396 2517 8397
rect 2451 8332 2452 8396
rect 2516 8332 2517 8396
rect 2451 8331 2517 8332
rect 2267 7308 2333 7309
rect 2267 7244 2268 7308
rect 2332 7244 2333 7308
rect 2267 7243 2333 7244
rect 2083 6900 2149 6901
rect 2083 6836 2084 6900
rect 2148 6836 2149 6900
rect 2083 6835 2149 6836
rect 1899 4044 1965 4045
rect 1899 3980 1900 4044
rect 1964 3980 1965 4044
rect 1899 3979 1965 3980
rect 1347 3092 1413 3093
rect 1347 3028 1348 3092
rect 1412 3028 1413 3092
rect 1347 3027 1413 3028
rect 1163 1596 1229 1597
rect 1163 1532 1164 1596
rect 1228 1532 1229 1596
rect 1163 1531 1229 1532
rect 2454 781 2514 8331
rect 2657 8192 2977 9216
rect 3187 9076 3253 9077
rect 3187 9012 3188 9076
rect 3252 9012 3253 9076
rect 3187 9011 3253 9012
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 3190 3365 3250 9011
rect 3371 6220 3437 6221
rect 3371 6156 3372 6220
rect 3436 6156 3437 6220
rect 3371 6155 3437 6156
rect 3187 3364 3253 3365
rect 3187 3300 3188 3364
rect 3252 3300 3253 3364
rect 3187 3299 3253 3300
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 3374 2685 3434 6155
rect 3558 3501 3618 9419
rect 3739 8940 3805 8941
rect 3739 8876 3740 8940
rect 3804 8876 3805 8940
rect 3739 8875 3805 8876
rect 3742 4181 3802 8875
rect 3926 7037 3986 12139
rect 3923 7036 3989 7037
rect 3923 6972 3924 7036
rect 3988 6972 3989 7036
rect 3923 6971 3989 6972
rect 3923 4588 3989 4589
rect 3923 4524 3924 4588
rect 3988 4524 3989 4588
rect 3923 4523 3989 4524
rect 3739 4180 3805 4181
rect 3739 4116 3740 4180
rect 3804 4116 3805 4180
rect 3739 4115 3805 4116
rect 3555 3500 3621 3501
rect 3555 3436 3556 3500
rect 3620 3436 3621 3500
rect 3555 3435 3621 3436
rect 3371 2684 3437 2685
rect 3371 2620 3372 2684
rect 3436 2620 3437 2684
rect 3371 2619 3437 2620
rect 3926 2549 3986 4523
rect 4110 2685 4170 12955
rect 4370 12000 4690 13024
rect 6084 16896 6404 17456
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 5579 13020 5645 13021
rect 5579 12956 5580 13020
rect 5644 12956 5645 13020
rect 5579 12955 5645 12956
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4843 10708 4909 10709
rect 4843 10644 4844 10708
rect 4908 10644 4909 10708
rect 4843 10643 4909 10644
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 3923 2548 3989 2549
rect 3923 2484 3924 2548
rect 3988 2484 3989 2548
rect 3923 2483 3989 2484
rect 4370 2208 4690 3232
rect 4846 2821 4906 10643
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5398 4045 5458 10235
rect 5582 4045 5642 12955
rect 5947 12612 6013 12613
rect 5947 12548 5948 12612
rect 6012 12548 6013 12612
rect 5947 12547 6013 12548
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 5579 4044 5645 4045
rect 5579 3980 5580 4044
rect 5644 3980 5645 4044
rect 5579 3979 5645 3980
rect 5950 3773 6010 12547
rect 6084 12544 6404 13568
rect 7797 17440 8117 17456
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 9511 16896 9831 17456
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 8339 14516 8405 14517
rect 8339 14452 8340 14516
rect 8404 14452 8405 14516
rect 8339 14451 8405 14452
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 6499 13156 6565 13157
rect 6499 13092 6500 13156
rect 6564 13092 6565 13156
rect 6499 13091 6565 13092
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6502 4045 6562 13091
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7419 12884 7485 12885
rect 7419 12820 7420 12884
rect 7484 12820 7485 12884
rect 7419 12819 7485 12820
rect 7051 12204 7117 12205
rect 7051 12140 7052 12204
rect 7116 12140 7117 12204
rect 7051 12139 7117 12140
rect 6867 9076 6933 9077
rect 6867 9012 6868 9076
rect 6932 9012 6933 9076
rect 6867 9011 6933 9012
rect 6683 7988 6749 7989
rect 6683 7924 6684 7988
rect 6748 7924 6749 7988
rect 6683 7923 6749 7924
rect 6686 4861 6746 7923
rect 6683 4860 6749 4861
rect 6683 4796 6684 4860
rect 6748 4796 6749 4860
rect 6683 4795 6749 4796
rect 6499 4044 6565 4045
rect 6499 3980 6500 4044
rect 6564 3980 6565 4044
rect 6499 3979 6565 3980
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 5947 3772 6013 3773
rect 5947 3708 5948 3772
rect 6012 3708 6013 3772
rect 5947 3707 6013 3708
rect 4843 2820 4909 2821
rect 4843 2756 4844 2820
rect 4908 2756 4909 2820
rect 4843 2755 4909 2756
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 2752 6404 3776
rect 6502 2821 6562 3979
rect 6870 3229 6930 9011
rect 6867 3228 6933 3229
rect 6867 3164 6868 3228
rect 6932 3164 6933 3228
rect 6867 3163 6933 3164
rect 7054 2821 7114 12139
rect 7422 3093 7482 12819
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 8342 6357 8402 14451
rect 8523 14380 8589 14381
rect 8523 14316 8524 14380
rect 8588 14316 8589 14380
rect 8523 14315 8589 14316
rect 8526 8261 8586 14315
rect 9075 13972 9141 13973
rect 9075 13908 9076 13972
rect 9140 13908 9141 13972
rect 9075 13907 9141 13908
rect 8523 8260 8589 8261
rect 8523 8196 8524 8260
rect 8588 8196 8589 8260
rect 8523 8195 8589 8196
rect 8339 6356 8405 6357
rect 8339 6292 8340 6356
rect 8404 6292 8405 6356
rect 8339 6291 8405 6292
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7419 3092 7485 3093
rect 7419 3028 7420 3092
rect 7484 3028 7485 3092
rect 7419 3027 7485 3028
rect 6499 2820 6565 2821
rect 6499 2756 6500 2820
rect 6564 2756 6565 2820
rect 6499 2755 6565 2756
rect 7051 2820 7117 2821
rect 7051 2756 7052 2820
rect 7116 2756 7117 2820
rect 7051 2755 7117 2756
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 2208 8117 3232
rect 9078 2549 9138 13907
rect 9511 13632 9831 14656
rect 11224 17440 11544 17456
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 9995 13836 10061 13837
rect 9995 13772 9996 13836
rect 10060 13772 10061 13836
rect 9995 13771 10061 13772
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9998 4725 10058 13771
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 12938 16896 13258 17456
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12571 11252 12637 11253
rect 12571 11188 12572 11252
rect 12636 11188 12637 11252
rect 12571 11187 12637 11188
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 10179 10572 10245 10573
rect 10179 10508 10180 10572
rect 10244 10508 10245 10572
rect 10179 10507 10245 10508
rect 9995 4724 10061 4725
rect 9995 4660 9996 4724
rect 10060 4660 10061 4724
rect 9995 4659 10061 4660
rect 9995 4316 10061 4317
rect 9995 4252 9996 4316
rect 10060 4252 10061 4316
rect 9995 4251 10061 4252
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9075 2548 9141 2549
rect 9075 2484 9076 2548
rect 9140 2484 9141 2548
rect 9075 2483 9141 2484
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 2128 9831 2688
rect 9998 1461 10058 4251
rect 10182 2277 10242 10507
rect 10363 10164 10429 10165
rect 10363 10100 10364 10164
rect 10428 10100 10429 10164
rect 10363 10099 10429 10100
rect 10366 9349 10426 10099
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 10363 9348 10429 9349
rect 10363 9284 10364 9348
rect 10428 9284 10429 9348
rect 10363 9283 10429 9284
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 10363 8532 10429 8533
rect 10363 8468 10364 8532
rect 10428 8468 10429 8532
rect 10363 8467 10429 8468
rect 10366 2685 10426 8467
rect 10731 7852 10797 7853
rect 10731 7788 10732 7852
rect 10796 7788 10797 7852
rect 10731 7787 10797 7788
rect 10734 2685 10794 7787
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 10915 7308 10981 7309
rect 10915 7244 10916 7308
rect 10980 7244 10981 7308
rect 10915 7243 10981 7244
rect 10918 4045 10978 7243
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 12574 6493 12634 11187
rect 12755 11116 12821 11117
rect 12755 11052 12756 11116
rect 12820 11052 12821 11116
rect 12755 11051 12821 11052
rect 12571 6492 12637 6493
rect 12571 6428 12572 6492
rect 12636 6428 12637 6492
rect 12571 6427 12637 6428
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 10915 4044 10981 4045
rect 10915 3980 10916 4044
rect 10980 3980 10981 4044
rect 10915 3979 10981 3980
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 10731 2684 10797 2685
rect 10731 2620 10732 2684
rect 10796 2620 10797 2684
rect 10731 2619 10797 2620
rect 10179 2276 10245 2277
rect 10179 2212 10180 2276
rect 10244 2212 10245 2276
rect 10179 2211 10245 2212
rect 11224 2208 11544 3232
rect 12758 2957 12818 11051
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12755 2956 12821 2957
rect 12755 2892 12756 2956
rect 12820 2892 12821 2956
rect 12755 2891 12821 2892
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 17440 14971 17456
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
rect 9995 1460 10061 1461
rect 9995 1396 9996 1460
rect 10060 1396 10061 1460
rect 9995 1395 10061 1396
rect 2451 780 2517 781
rect 2451 716 2452 780
rect 2516 716 2517 780
rect 2451 715 2517 716
use sky130_fd_sc_hd__inv_2  _177_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _178_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _180_
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _184_
timestamp 1688980957
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _185_
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _191_
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1688980957
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _193_
timestamp 1688980957
transform 1 0 13248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1688980957
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1688980957
transform 1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1688980957
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1688980957
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1688980957
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform 1 0 10580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1688980957
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1688980957
transform 1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1688980957
transform 1 0 5336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _231_
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _232_
timestamp 1688980957
transform 1 0 3036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1688980957
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1688980957
transform 1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _235_
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1688980957
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1688980957
transform 1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1688980957
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1688980957
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform 1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform 1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1688980957
transform 1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _254_
timestamp 1688980957
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1688980957
transform 1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1688980957
transform 1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1688980957
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1688980957
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1688980957
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1688980957
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1688980957
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1688980957
transform 1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1688980957
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1688980957
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1688980957
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1688980957
transform 1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1688980957
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1688980957
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1688980957
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _293_
timestamp 1688980957
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _295_
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1688980957
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1688980957
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1688980957
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1688980957
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1688980957
transform 1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1688980957
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1688980957
transform 1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1688980957
transform 1 0 13248 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1688980957
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1688980957
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1688980957
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1688980957
transform 1 0 11592 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1688980957
transform 1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1688980957
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1688980957
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1688980957
transform 1 0 5612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1688980957
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1688980957
transform 1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1688980957
transform 1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1688980957
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1688980957
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1688980957
transform 1 0 1472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1688980957
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1688980957
transform 1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1688980957
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1688980957
transform 1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1688980957
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1688980957
transform 1 0 9108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1688980957
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1688980957
transform 1 0 8464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1688980957
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1688980957
transform 1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _387_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1688980957
transform 1 0 10488 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _389_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1688980957
transform 1 0 4692 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _392_
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _395_
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1688980957
transform 1 0 1472 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _398_
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _406_
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _421_
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _422_
timestamp 1688980957
transform 1 0 9292 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _439_
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _440_
timestamp 1688980957
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _441_
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _442_
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _443_
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _445_
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _447_
timestamp 1688980957
transform 1 0 12144 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _449_
timestamp 1688980957
transform 1 0 12420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _450_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _451_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _452_
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _453_
timestamp 1688980957
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _454_
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _455_
timestamp 1688980957
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _455__63 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _456_
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _457_
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _458_
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _459_
timestamp 1688980957
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _460_
timestamp 1688980957
transform 1 0 10764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _461_
timestamp 1688980957
transform 1 0 12788 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _462_
timestamp 1688980957
transform 1 0 6992 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _463__64
timestamp 1688980957
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _463_
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _464_
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _465_
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _466_
timestamp 1688980957
transform 1 0 3956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _467_
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _468_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _469_
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _470_
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _471_
timestamp 1688980957
transform 1 0 6624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _472_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _473_
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _474_
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _475__65
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _475_
timestamp 1688980957
transform 1 0 1840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _476_
timestamp 1688980957
transform 1 0 4416 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _477_
timestamp 1688980957
transform 1 0 1840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _478_
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _479_
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _480_
timestamp 1688980957
transform 1 0 2944 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _481_
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _482_
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _483_
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _484_
timestamp 1688980957
transform 1 0 3036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _485_
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _486_
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _487__66
timestamp 1688980957
transform 1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _487_
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _488_
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _489_
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _490_
timestamp 1688980957
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _491_
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _492_
timestamp 1688980957
transform 1 0 4048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _493_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _494_
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _495_
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _496_
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _497_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _498_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _499__67
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _499_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _500_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _501_
timestamp 1688980957
transform 1 0 5152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _502_
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _503_
timestamp 1688980957
transform 1 0 5704 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _504_
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _505_
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _506_
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _507_
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _508_
timestamp 1688980957
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _509__68
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _509_
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _510_
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _511_
timestamp 1688980957
transform 1 0 7636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _512_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _513_
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _514_
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _515_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _516_
timestamp 1688980957
transform 1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _517_
timestamp 1688980957
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _518_
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _519__69
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _519_
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _520_
timestamp 1688980957
transform 1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _521_
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _522_
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _523_
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _524_
timestamp 1688980957
transform 1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _525_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _525__70
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _526_
timestamp 1688980957
transform 1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _527_
timestamp 1688980957
transform 1 0 8004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _528_
timestamp 1688980957
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _529_
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _530__71
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _530_
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _531_
timestamp 1688980957
transform 1 0 9752 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _532_
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _533_
timestamp 1688980957
transform 1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _534__72
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _534_
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _535_
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _536_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _537_
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _538__73
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _538_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _539_
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _540_
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _541_
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _542_
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _542__74
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _543_
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _544_
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _545_
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _546__75
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _546_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _547_
timestamp 1688980957
transform 1 0 13248 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _548_
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _549_
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _550_
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _550__76
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _551_
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _552_
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _553_
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _554__77
timestamp 1688980957
transform 1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _554_
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _555_
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _556_
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _557_
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 1564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 1840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_prog_clk
timestamp 1688980957
transform 1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_prog_clk
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_19
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_38
timestamp 1688980957
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_94
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_16
timestamp 1688980957
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_88
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_116
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_144
timestamp 1688980957
transform 1 0 14352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_20
timestamp 1688980957
transform 1 0 2944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_37
timestamp 1688980957
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_91
timestamp 1688980957
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_32
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_104
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_108
timestamp 1688980957
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_52
timestamp 1688980957
transform 1 0 5888 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_71
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_99
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_19
timestamp 1688980957
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_49
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_79
timestamp 1688980957
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_45
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_67
timestamp 1688980957
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_108
timestamp 1688980957
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_118
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_144
timestamp 1688980957
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_144
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_144
timestamp 1688980957
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_8
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_17
timestamp 1688980957
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_91
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_10
timestamp 1688980957
transform 1 0 2024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_135
timestamp 1688980957
transform 1 0 13524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_20
timestamp 1688980957
transform 1 0 2944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_6
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_10
timestamp 1688980957
transform 1 0 2024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_28
timestamp 1688980957
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_77
timestamp 1688980957
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_12
timestamp 1688980957
transform 1 0 2208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_55
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_101
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_144
timestamp 1688980957
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_6
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_79 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_91
timestamp 1688980957
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_95
timestamp 1688980957
transform 1 0 9844 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1688980957
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_127
timestamp 1688980957
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_96
timestamp 1688980957
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_20
timestamp 1688980957
transform 1 0 2944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_24
timestamp 1688980957
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_124
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_144
timestamp 1688980957
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_17
timestamp 1688980957
transform 1 0 2668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_39
timestamp 1688980957
transform 1 0 4692 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_46
timestamp 1688980957
transform 1 0 5336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_135
timestamp 1688980957
transform 1 0 13524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_37
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_41
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_73
timestamp 1688980957
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_90
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_103
timestamp 1688980957
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_128
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_16
timestamp 1688980957
transform 1 0 2576 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_20
timestamp 1688980957
transform 1 0 2944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_33
timestamp 1688980957
transform 1 0 4140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_45
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_69
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_88
timestamp 1688980957
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_105
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_117
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_129
timestamp 1688980957
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_6
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_10
timestamp 1688980957
transform 1 0 2024 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_36
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp 1688980957
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_52
timestamp 1688980957
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_64
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_21
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_45
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_145
timestamp 1688980957
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_14
timestamp 1688980957
transform 1 0 2392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_80
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_19
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 12696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 10764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 8740 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 12696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 13524 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 7728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 11960 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 6532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 1564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 6624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 2668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 14260 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform 1 0 2300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1688980957
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1688980957
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1688980957
transform 1 0 14168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output54
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1688980957
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output57
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 0 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
flabel metal3 s 15200 17688 16000 17808 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 15200 18504 16000 18624 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 5 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 6 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 7 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 8 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 9 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 10 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 11 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 12 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 13 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 14 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 15 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 16 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 17 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 18 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 19 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 20 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 21 nsew signal tristate
flabel metal3 s 15200 1368 16000 1488 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 22 nsew signal input
flabel metal3 s 15200 2184 16000 2304 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 23 nsew signal input
flabel metal3 s 15200 3000 16000 3120 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 24 nsew signal input
flabel metal3 s 15200 3816 16000 3936 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 25 nsew signal input
flabel metal3 s 15200 4632 16000 4752 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 26 nsew signal input
flabel metal3 s 15200 5448 16000 5568 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 27 nsew signal input
flabel metal3 s 15200 6264 16000 6384 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 28 nsew signal input
flabel metal3 s 15200 7080 16000 7200 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 29 nsew signal input
flabel metal3 s 15200 7896 16000 8016 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 30 nsew signal input
flabel metal3 s 15200 8712 16000 8832 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal3 s 15200 9528 16000 9648 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 32 nsew signal tristate
flabel metal3 s 15200 10344 16000 10464 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 33 nsew signal tristate
flabel metal3 s 15200 11160 16000 11280 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 34 nsew signal tristate
flabel metal3 s 15200 11976 16000 12096 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 35 nsew signal tristate
flabel metal3 s 15200 12792 16000 12912 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 36 nsew signal tristate
flabel metal3 s 15200 13608 16000 13728 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 37 nsew signal tristate
flabel metal3 s 15200 14424 16000 14544 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 38 nsew signal tristate
flabel metal3 s 15200 15240 16000 15360 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 39 nsew signal tristate
flabel metal2 s 570 0 626 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 40 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 41 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 42 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 43 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 44 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 45 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 46 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 47 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 48 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 49 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 50 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 51 nsew signal tristate
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 52 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 53 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 54 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 55 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 56 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 57 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 58 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 59 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 prog_clk
port 60 nsew signal input
flabel metal3 s 15200 16056 16000 16176 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 61 nsew signal input
flabel metal3 s 15200 16872 16000 16992 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 62 nsew signal input
flabel metal4 s 2657 2128 2977 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 6084 2128 6404 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 9511 2128 9831 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 12938 2128 13258 17456 0 FreeSans 1920 90 0 0 vdd
port 63 nsew power bidirectional
flabel metal4 s 4370 2128 4690 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 17456 0 FreeSans 1920 90 0 0 vss
port 64 nsew ground bidirectional
rlabel metal1 7958 16864 7958 16864 0 vdd
rlabel via1 8037 17408 8037 17408 0 vss
rlabel metal1 2438 2040 2438 2040 0 _000_
rlabel metal1 1472 3706 1472 3706 0 _001_
rlabel metal1 6716 5338 6716 5338 0 _002_
rlabel metal1 11592 3706 11592 3706 0 _003_
rlabel metal1 13018 12784 13018 12784 0 _004_
rlabel metal1 13340 12818 13340 12818 0 _005_
rlabel metal1 14490 5236 14490 5236 0 _006_
rlabel metal1 13524 8942 13524 8942 0 _007_
rlabel via2 11730 6307 11730 6307 0 _008_
rlabel metal1 14214 2618 14214 2618 0 _009_
rlabel metal1 7912 7242 7912 7242 0 _010_
rlabel metal1 9246 6324 9246 6324 0 _011_
rlabel metal1 9936 9554 9936 9554 0 _012_
rlabel metal1 9844 8602 9844 8602 0 _013_
rlabel metal1 4462 3706 4462 3706 0 _014_
rlabel metal1 9292 3162 9292 3162 0 _015_
rlabel metal1 7682 4148 7682 4148 0 _016_
rlabel metal1 5934 4250 5934 4250 0 _017_
rlabel metal1 7079 9418 7079 9418 0 _018_
rlabel metal2 2162 13124 2162 13124 0 _019_
rlabel metal1 8326 11152 8326 11152 0 _020_
rlabel metal1 9522 12852 9522 12852 0 _021_
rlabel metal1 7360 11866 7360 11866 0 _022_
rlabel metal1 10488 14382 10488 14382 0 _023_
rlabel metal1 7866 13430 7866 13430 0 _024_
rlabel metal1 2576 12410 2576 12410 0 _025_
rlabel metal1 4140 13838 4140 13838 0 _026_
rlabel metal2 1058 8177 1058 8177 0 _027_
rlabel metal1 6256 5066 6256 5066 0 _028_
rlabel metal1 3588 5882 3588 5882 0 _029_
rlabel metal1 5750 6188 5750 6188 0 _030_
rlabel metal1 2599 7990 2599 7990 0 _031_
rlabel metal1 1702 5882 1702 5882 0 _032_
rlabel metal1 4416 11730 4416 11730 0 _033_
rlabel metal1 1886 9690 1886 9690 0 _034_
rlabel metal2 3450 11560 3450 11560 0 _035_
rlabel metal1 13202 4046 13202 4046 0 _036_
rlabel metal2 3266 11356 3266 11356 0 _037_
rlabel metal1 3450 14416 3450 14416 0 _038_
rlabel metal2 3404 12614 3404 12614 0 _039_
rlabel metal2 1794 8908 1794 8908 0 _040_
rlabel metal1 1472 11322 1472 11322 0 _041_
rlabel metal1 2300 9146 2300 9146 0 _042_
rlabel metal1 5474 9418 5474 9418 0 _043_
rlabel metal1 3910 9520 3910 9520 0 _044_
rlabel metal1 5658 10778 5658 10778 0 _045_
rlabel metal1 6348 8602 6348 8602 0 _046_
rlabel metal1 6118 9690 6118 9690 0 _047_
rlabel metal1 11362 12784 11362 12784 0 _048_
rlabel metal1 12466 11696 12466 11696 0 _049_
rlabel metal2 10166 12172 10166 12172 0 _050_
rlabel metal2 14214 10115 14214 10115 0 _051_
rlabel metal1 10718 10064 10718 10064 0 _052_
rlabel metal2 14306 11322 14306 11322 0 _053_
rlabel metal2 12466 12444 12466 12444 0 _054_
rlabel metal1 13938 10744 13938 10744 0 _055_
rlabel metal1 10120 11866 10120 11866 0 _056_
rlabel metal1 10718 10234 10718 10234 0 _057_
rlabel metal2 13202 12036 13202 12036 0 _058_
rlabel metal1 13524 10098 13524 10098 0 _059_
rlabel metal2 11730 9860 11730 9860 0 _060_
rlabel metal1 12926 11730 12926 11730 0 _061_
rlabel metal1 12650 10098 12650 10098 0 _062_
rlabel metal2 13386 10336 13386 10336 0 _063_
rlabel metal1 10672 11866 10672 11866 0 _064_
rlabel metal2 13018 13124 13018 13124 0 _065_
rlabel metal1 7222 11016 7222 11016 0 _066_
rlabel metal1 6716 11118 6716 11118 0 _067_
rlabel metal1 6394 9486 6394 9486 0 _068_
rlabel metal1 6854 9044 6854 9044 0 _069_
rlabel metal1 4186 9452 4186 9452 0 _070_
rlabel metal1 2714 9452 2714 9452 0 _071_
rlabel metal1 6854 10166 6854 10166 0 _072_
rlabel metal1 7084 10234 7084 10234 0 _073_
rlabel metal1 5290 9554 5290 9554 0 _074_
rlabel metal1 6854 8500 6854 8500 0 _075_
rlabel metal1 3772 9010 3772 9010 0 _076_
rlabel metal2 5750 9588 5750 9588 0 _077_
rlabel metal2 3588 12172 3588 12172 0 _078_
rlabel metal3 1863 12580 1863 12580 0 _079_
rlabel metal1 4784 4590 4784 4590 0 _080_
rlabel metal1 1978 3570 1978 3570 0 _081_
rlabel metal1 1518 3366 1518 3366 0 _082_
rlabel metal1 12834 3910 12834 3910 0 _083_
rlabel metal2 2438 6800 2438 6800 0 _084_
rlabel metal1 2346 4760 2346 4760 0 _085_
rlabel metal1 3680 4046 3680 4046 0 _086_
rlabel via2 2438 4029 2438 4029 0 _087_
rlabel metal3 1679 13804 1679 13804 0 _088_
rlabel metal1 3772 3162 3772 3162 0 _089_
rlabel metal1 4140 12886 4140 12886 0 _090_
rlabel metal2 2898 12002 2898 12002 0 _091_
rlabel metal1 2898 8058 2898 8058 0 _092_
rlabel metal1 2346 10540 2346 10540 0 _093_
rlabel metal1 2392 7242 2392 7242 0 _094_
rlabel metal2 5474 7412 5474 7412 0 _095_
rlabel metal1 4646 12886 4646 12886 0 _096_
rlabel metal1 3634 11186 3634 11186 0 _097_
rlabel metal1 3174 7956 3174 7956 0 _098_
rlabel metal1 3588 10098 3588 10098 0 _099_
rlabel metal1 2070 7514 2070 7514 0 _100_
rlabel metal2 7314 7650 7314 7650 0 _101_
rlabel metal2 4830 6052 4830 6052 0 _102_
rlabel metal1 3956 6426 3956 6426 0 _103_
rlabel metal1 5750 13838 5750 13838 0 _104_
rlabel metal2 1978 4233 1978 4233 0 _105_
rlabel metal2 1242 13231 1242 13231 0 _106_
rlabel metal1 4968 5882 4968 5882 0 _107_
rlabel metal1 4646 7412 4646 7412 0 _108_
rlabel metal2 1794 4658 1794 4658 0 _109_
rlabel metal1 10097 4726 10097 4726 0 _110_
rlabel metal1 1472 2618 1472 2618 0 _111_
rlabel metal1 9614 14280 9614 14280 0 _112_
rlabel metal1 8280 13362 8280 13362 0 _113_
rlabel metal1 9062 12750 9062 12750 0 _114_
rlabel metal1 7866 12342 7866 12342 0 _115_
rlabel metal1 9154 11220 9154 11220 0 _116_
rlabel metal1 10074 13974 10074 13974 0 _117_
rlabel metal1 7958 13498 7958 13498 0 _118_
rlabel metal1 9476 12274 9476 12274 0 _119_
rlabel metal1 8188 11730 8188 11730 0 _120_
rlabel metal1 8694 10642 8694 10642 0 _121_
rlabel metal4 1196 7888 1196 7888 0 _122_
rlabel metal3 1587 10812 1587 10812 0 _123_
rlabel metal1 7130 5338 7130 5338 0 _124_
rlabel metal1 7130 3094 7130 3094 0 _125_
rlabel metal1 1564 13362 1564 13362 0 _126_
rlabel metal1 6256 2958 6256 2958 0 _127_
rlabel metal1 8878 3128 8878 3128 0 _128_
rlabel metal2 7498 4352 7498 4352 0 _129_
rlabel metal1 5520 4658 5520 4658 0 _130_
rlabel metal1 8418 3434 8418 3434 0 _131_
rlabel metal1 8464 4114 8464 4114 0 _132_
rlabel metal2 2990 2040 2990 2040 0 _133_
rlabel metal1 10304 8534 10304 8534 0 _134_
rlabel metal1 9614 9690 9614 9690 0 _135_
rlabel metal2 10626 9112 10626 9112 0 _136_
rlabel metal1 9476 10166 9476 10166 0 _137_
rlabel metal1 9522 6392 9522 6392 0 _138_
rlabel metal1 8142 7922 8142 7922 0 _139_
rlabel metal1 9154 6664 9154 6664 0 _140_
rlabel metal1 7958 5882 7958 5882 0 _141_
rlabel metal1 13800 5882 13800 5882 0 _142_
rlabel metal1 10810 5746 10810 5746 0 _143_
rlabel metal1 10166 2618 10166 2618 0 _144_
rlabel metal1 11224 5746 11224 5746 0 _145_
rlabel metal1 13340 7786 13340 7786 0 _146_
rlabel metal1 14260 5338 14260 5338 0 _147_
rlabel metal2 14398 7480 14398 7480 0 _148_
rlabel metal1 14168 8058 14168 8058 0 _149_
rlabel metal1 13524 12614 13524 12614 0 _150_
rlabel metal1 13248 12614 13248 12614 0 _151_
rlabel metal1 14398 12614 14398 12614 0 _152_
rlabel metal1 13570 7446 13570 7446 0 _153_
rlabel metal2 11776 2346 11776 2346 0 _154_
rlabel metal1 10856 2482 10856 2482 0 _155_
rlabel metal1 13386 2312 13386 2312 0 _156_
rlabel via2 1518 2907 1518 2907 0 _157_
rlabel metal2 12558 5185 12558 5185 0 _158_
rlabel metal2 4002 2006 4002 2006 0 _159_
rlabel metal2 11822 12019 11822 12019 0 _160_
rlabel metal1 4784 2618 4784 2618 0 _161_
rlabel metal2 7958 823 7958 823 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 7222 823 7222 823 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 14536 17170 14536 17170 0 ccff_head
rlabel metal1 13800 17306 13800 17306 0 ccff_tail
rlabel metal3 1027 3060 1027 3060 0 chanx_left_in[0]
rlabel metal3 1027 3876 1027 3876 0 chanx_left_in[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_in[2]
rlabel metal3 1188 5508 1188 5508 0 chanx_left_in[3]
rlabel metal3 1050 6324 1050 6324 0 chanx_left_in[4]
rlabel metal3 1027 7140 1027 7140 0 chanx_left_in[5]
rlabel metal3 1027 7956 1027 7956 0 chanx_left_in[6]
rlabel metal3 843 8772 843 8772 0 chanx_left_in[7]
rlabel metal3 820 9588 820 9588 0 chanx_left_in[8]
rlabel metal3 820 12036 820 12036 0 chanx_left_out[0]
rlabel metal3 820 12852 820 12852 0 chanx_left_out[1]
rlabel metal3 1142 13668 1142 13668 0 chanx_left_out[2]
rlabel metal3 820 14484 820 14484 0 chanx_left_out[3]
rlabel metal3 912 15300 912 15300 0 chanx_left_out[4]
rlabel metal3 820 16116 820 16116 0 chanx_left_out[5]
rlabel metal3 866 16932 866 16932 0 chanx_left_out[6]
rlabel metal3 820 17748 820 17748 0 chanx_left_out[7]
rlabel metal2 2806 17901 2806 17901 0 chanx_left_out[8]
rlabel metal2 8096 2346 8096 2346 0 chanx_right_in[0]
rlabel metal1 3082 14382 3082 14382 0 chanx_right_in[1]
rlabel metal1 14076 3026 14076 3026 0 chanx_right_in[2]
rlabel metal2 8418 3672 8418 3672 0 chanx_right_in[3]
rlabel metal1 13938 3502 13938 3502 0 chanx_right_in[4]
rlabel metal2 2622 2465 2622 2465 0 chanx_right_in[5]
rlabel metal1 13754 13260 13754 13260 0 chanx_right_in[6]
rlabel metal2 13754 8041 13754 8041 0 chanx_right_in[7]
rlabel metal3 3289 2652 3289 2652 0 chanx_right_in[8]
rlabel metal2 14398 8993 14398 8993 0 chanx_right_out[0]
rlabel via2 14122 9571 14122 9571 0 chanx_right_out[1]
rlabel metal2 14398 10319 14398 10319 0 chanx_right_out[2]
rlabel metal2 14398 11373 14398 11373 0 chanx_right_out[3]
rlabel metal2 14398 12257 14398 12257 0 chanx_right_out[4]
rlabel metal2 14398 13005 14398 13005 0 chanx_right_out[5]
rlabel metal1 14444 13838 14444 13838 0 chanx_right_out[6]
rlabel metal2 14398 14637 14398 14637 0 chanx_right_out[7]
rlabel metal1 14628 15674 14628 15674 0 chanx_right_out[8]
rlabel metal1 1288 2958 1288 2958 0 chany_bottom_in[0]
rlabel metal2 1334 823 1334 823 0 chany_bottom_in[1]
rlabel metal2 2208 5372 2208 5372 0 chany_bottom_in[2]
rlabel metal2 2806 823 2806 823 0 chany_bottom_in[3]
rlabel metal2 3542 1826 3542 1826 0 chany_bottom_in[4]
rlabel metal1 1794 14246 1794 14246 0 chany_bottom_in[5]
rlabel metal2 5014 1044 5014 1044 0 chany_bottom_in[6]
rlabel metal1 9246 13736 9246 13736 0 chany_bottom_in[7]
rlabel metal2 6486 823 6486 823 0 chany_bottom_in[8]
rlabel metal2 8694 1520 8694 1520 0 chany_bottom_out[0]
rlabel metal2 9430 1554 9430 1554 0 chany_bottom_out[1]
rlabel metal2 10166 1792 10166 1792 0 chany_bottom_out[2]
rlabel metal1 12650 5576 12650 5576 0 chany_bottom_out[3]
rlabel metal2 13846 3672 13846 3672 0 chany_bottom_out[4]
rlabel metal1 8510 2414 8510 2414 0 chany_bottom_out[5]
rlabel metal2 13110 1418 13110 1418 0 chany_bottom_out[6]
rlabel metal2 13846 823 13846 823 0 chany_bottom_out[7]
rlabel metal1 14214 3434 14214 3434 0 chany_bottom_out[8]
rlabel metal1 8050 7446 8050 7446 0 clknet_0_prog_clk
rlabel metal1 1426 6324 1426 6324 0 clknet_2_0__leaf_prog_clk
rlabel metal1 1518 10166 1518 10166 0 clknet_2_1__leaf_prog_clk
rlabel metal1 7912 4590 7912 4590 0 clknet_2_2__leaf_prog_clk
rlabel metal1 10120 13294 10120 13294 0 clknet_2_3__leaf_prog_clk
rlabel metal3 820 10404 820 10404 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 2116 14994 2116 14994 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 6716 6222 6716 6222 0 mem_bottom_track_1.DFF_0_.D
rlabel metal1 6624 5882 6624 5882 0 mem_bottom_track_1.DFF_0_.Q
rlabel viali 5377 8942 5377 8942 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal1 9798 2414 9798 2414 0 mem_bottom_track_11.DFF_0_.D
rlabel metal2 12926 8772 12926 8772 0 mem_bottom_track_11.DFF_0_.Q
rlabel metal1 12788 7310 12788 7310 0 mem_bottom_track_11.DFF_1_.Q
rlabel metal1 14260 12750 14260 12750 0 mem_bottom_track_13.DFF_0_.Q
rlabel metal1 13846 12818 13846 12818 0 mem_bottom_track_13.DFF_1_.Q
rlabel metal1 6394 5202 6394 5202 0 mem_bottom_track_15.DFF_0_.Q
rlabel metal1 11684 3502 11684 3502 0 mem_bottom_track_15.DFF_1_.Q
rlabel metal1 4462 2414 4462 2414 0 mem_bottom_track_17.DFF_0_.Q
rlabel metal3 5865 12580 5865 12580 0 mem_bottom_track_17.DFF_1_.Q
rlabel metal1 4830 3468 4830 3468 0 mem_bottom_track_3.DFF_0_.Q
rlabel metal1 9706 3060 9706 3060 0 mem_bottom_track_3.DFF_1_.Q
rlabel metal1 10212 6222 10212 6222 0 mem_bottom_track_5.DFF_0_.Q
rlabel metal1 10074 9452 10074 9452 0 mem_bottom_track_5.DFF_1_.Q
rlabel metal2 7682 8330 7682 8330 0 mem_bottom_track_7.DFF_0_.Q
rlabel metal1 10212 6766 10212 6766 0 mem_bottom_track_7.DFF_1_.Q
rlabel metal1 10534 7174 10534 7174 0 mem_bottom_track_9.DFF_0_.Q
rlabel metal1 2254 13940 2254 13940 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 2162 11220 2162 11220 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 3220 10574 3220 10574 0 mem_left_track_1.DFF_2_.Q
rlabel metal2 4646 12619 4646 12619 0 mem_left_track_17.DFF_0_.D
rlabel metal1 6762 12206 6762 12206 0 mem_left_track_17.DFF_0_.Q
rlabel metal1 8602 12818 8602 12818 0 mem_left_track_17.DFF_1_.Q
rlabel metal2 5980 6290 5980 6290 0 mem_left_track_9.DFF_0_.Q
rlabel metal1 2898 9928 2898 9928 0 mem_left_track_9.DFF_1_.Q
rlabel metal2 11224 9554 11224 9554 0 mem_right_track_0.DFF_0_.Q
rlabel metal1 12558 11764 12558 11764 0 mem_right_track_0.DFF_1_.Q
rlabel metal1 13386 9554 13386 9554 0 mem_right_track_0.DFF_2_.Q
rlabel metal1 5382 9996 5382 9996 0 mem_right_track_16.DFF_0_.D
rlabel metal1 10442 4556 10442 4556 0 mem_right_track_16.DFF_0_.Q
rlabel metal1 3634 5712 3634 5712 0 mem_right_track_16.DFF_1_.Q
rlabel metal1 6716 9554 6716 9554 0 mem_right_track_8.DFF_0_.Q
rlabel metal1 5382 9622 5382 9622 0 mem_right_track_8.DFF_1_.Q
rlabel metal1 3542 2584 3542 2584 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 6394 7174 6394 7174 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal2 4830 3468 4830 3468 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 7314 2958 7314 2958 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 6302 2482 6302 2482 0 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 4416 13974 4416 13974 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11500 9078 11500 9078 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal1 12650 9384 12650 9384 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal1 12880 8534 12880 8534 0 mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13662 7786 13662 7786 0 mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13386 7276 13386 7276 0 mux_bottom_track_13.INVTX1_0_.out
rlabel metal1 9338 4114 9338 4114 0 mux_bottom_track_13.INVTX1_1_.out
rlabel metal1 13294 5780 13294 5780 0 mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14260 5066 14260 5066 0 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5336 3366 5336 3366 0 mux_bottom_track_15.INVTX1_0_.out
rlabel metal2 10442 4641 10442 4641 0 mux_bottom_track_15.INVTX1_1_.out
rlabel metal2 12834 2550 12834 2550 0 mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13846 2584 13846 2584 0 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 12006 7548 12006 7548 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 3542 13940 3542 13940 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 12512 5542 12512 5542 0 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13202 2550 13202 2550 0 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal3 6325 12852 6325 12852 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal1 5152 4590 5152 4590 0 mux_bottom_track_3.INVTX1_1_.out
rlabel via2 1518 7803 1518 7803 0 mux_bottom_track_3.INVTX1_2_.out
rlabel metal1 8142 3604 8142 3604 0 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9108 4250 9108 4250 0 mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 6624 2006 6624 2006 0 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8924 11118 8924 11118 0 mux_bottom_track_5.INVTX1_0_.out
rlabel metal1 10120 10574 10120 10574 0 mux_bottom_track_5.INVTX1_1_.out
rlabel metal1 10120 10234 10120 10234 0 mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4324 2278 4324 2278 0 mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7130 6222 7130 6222 0 mux_bottom_track_7.INVTX1_0_.out
rlabel metal2 6670 8466 6670 8466 0 mux_bottom_track_7.INVTX1_1_.out
rlabel metal1 8418 6426 8418 6426 0 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 7728 12614 7728 12614 0 mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 11316 5678 11316 5678 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 6113 8058 6113 8058 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal2 11638 6358 11638 6358 0 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 11822 6698 11822 6698 0 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 3312 4114 3312 4114 0 mux_left_track_1.INVTX1_2_.out
rlabel via2 2438 14467 2438 14467 0 mux_left_track_1.INVTX1_3_.out
rlabel metal3 5543 10268 5543 10268 0 mux_left_track_1.INVTX1_4_.out
rlabel metal4 2300 8568 2300 8568 0 mux_left_track_1.INVTX1_5_.out
rlabel metal1 10258 5134 10258 5134 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 3726 4386 3726 4386 0 mux_left_track_1.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 2530 3808 2530 3808 0 mux_left_track_1.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 4554 4794 4554 4794 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 2622 5610 2622 5610 0 mux_left_track_1.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 2070 11679 2070 11679 0 mux_left_track_1.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 9430 11662 9430 11662 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 10350 12274 10350 12274 0 mux_left_track_17.INVTX1_3_.out
rlabel metal2 4738 2108 4738 2108 0 mux_left_track_17.INVTX1_4_.out
rlabel metal1 9154 11322 9154 11322 0 mux_left_track_17.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 8464 12750 8464 12750 0 mux_left_track_17.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 9246 13328 9246 13328 0 mux_left_track_17.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9062 14042 9062 14042 0 mux_left_track_17.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 2162 16592 2162 16592 0 mux_left_track_17.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 1840 8398 1840 8398 0 mux_left_track_9.INVTX1_2_.out
rlabel metal1 2714 8908 2714 8908 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 4002 9588 4002 9588 0 mux_left_track_9.INVTX1_4_.out
rlabel metal1 1656 9690 1656 9690 0 mux_left_track_9.INVTX1_5_.out
rlabel metal1 4508 7786 4508 7786 0 mux_left_track_9.mux_l1_in_0_.TGATE_0_.out
rlabel via1 2714 8468 2714 8468 0 mux_left_track_9.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 3910 11118 3910 11118 0 mux_left_track_9.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 4186 10370 4186 10370 0 mux_left_track_9.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 3634 11662 3634 11662 0 mux_left_track_9.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 4186 13838 4186 13838 0 mux_left_track_9.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 12788 13362 12788 13362 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 13202 12410 13202 12410 0 mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 13018 12308 13018 12308 0 mux_right_track_0.mux_l1_in_1_.TGATE_0_.out
rlabel metal1 11638 10234 11638 10234 0 mux_right_track_0.mux_l1_in_2_.TGATE_0_.out
rlabel metal2 13662 11968 13662 11968 0 mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 13202 10166 13202 10166 0 mux_right_track_0.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 13708 11050 13708 11050 0 mux_right_track_0.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 4278 3638 4278 3638 0 mux_right_track_16.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 5566 4998 5566 4998 0 mux_right_track_16.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 5106 5491 5106 5491 0 mux_right_track_16.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5336 7242 5336 7242 0 mux_right_track_16.mux_l2_in_1_.TGATE_0_.out
rlabel metal1 7038 7208 7038 7208 0 mux_right_track_16.mux_l3_in_0_.TGATE_0_.out
rlabel metal2 5980 10098 5980 10098 0 mux_right_track_8.INVTX1_0_.out
rlabel metal1 6348 9894 6348 9894 0 mux_right_track_8.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 4462 9690 4462 9690 0 mux_right_track_8.mux_l1_in_1_.TGATE_0_.out
rlabel metal2 7222 9860 7222 9860 0 mux_right_track_8.mux_l1_in_2_.TGATE_0_.out
rlabel metal1 6118 9622 6118 9622 0 mux_right_track_8.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 7038 11050 7038 11050 0 mux_right_track_8.mux_l2_in_1_.TGATE_0_.out
rlabel metal2 13294 11526 13294 11526 0 mux_right_track_8.mux_l3_in_0_.TGATE_0_.out
rlabel metal1 5106 13328 5106 13328 0 net1
rlabel metal1 4508 14042 4508 14042 0 net10
rlabel metal2 8418 4386 8418 4386 0 net100
rlabel metal2 2162 9282 2162 9282 0 net101
rlabel via1 4089 6766 4089 6766 0 net102
rlabel metal1 4595 10642 4595 10642 0 net103
rlabel metal2 12650 10846 12650 10846 0 net104
rlabel metal1 4921 6358 4921 6358 0 net105
rlabel metal1 2116 5338 2116 5338 0 net106
rlabel metal1 7171 12818 7171 12818 0 net107
rlabel metal1 5377 11050 5377 11050 0 net108
rlabel metal1 11495 11050 11495 11050 0 net109
rlabel metal1 1518 4114 1518 4114 0 net11
rlabel metal1 3082 11322 3082 11322 0 net110
rlabel metal1 5515 3434 5515 3434 0 net111
rlabel metal2 7038 4386 7038 4386 0 net112
rlabel metal2 1426 8330 1426 8330 0 net12
rlabel metal1 2760 3502 2760 3502 0 net13
rlabel metal1 8510 9520 8510 9520 0 net14
rlabel metal1 13018 9996 13018 9996 0 net15
rlabel metal1 3312 3162 3312 3162 0 net16
rlabel metal1 14214 3706 14214 3706 0 net17
rlabel metal1 6026 6188 6026 6188 0 net18
rlabel metal1 8602 16558 8602 16558 0 net19
rlabel metal1 2300 2414 2300 2414 0 net2
rlabel metal2 13570 8721 13570 8721 0 net20
rlabel metal2 3358 2329 3358 2329 0 net21
rlabel metal1 2254 3162 2254 3162 0 net22
rlabel metal1 2576 12614 2576 12614 0 net23
rlabel metal2 4278 7242 4278 7242 0 net24
rlabel metal1 2300 7854 2300 7854 0 net25
rlabel metal1 2530 15062 2530 15062 0 net26
rlabel metal1 2346 14416 2346 14416 0 net27
rlabel metal1 1978 12818 1978 12818 0 net28
rlabel metal3 4393 2652 4393 2652 0 net29
rlabel metal1 14306 13464 14306 13464 0 net3
rlabel metal1 5060 13226 5060 13226 0 net30
rlabel metal1 1472 9554 1472 9554 0 net31
rlabel metal2 3634 14331 3634 14331 0 net32
rlabel metal2 13846 16048 13846 16048 0 net33
rlabel metal1 13202 13906 13202 13906 0 net34
rlabel metal1 10856 14382 10856 14382 0 net35
rlabel metal1 1840 11866 1840 11866 0 net36
rlabel metal1 2162 2516 2162 2516 0 net37
rlabel metal2 1518 14161 1518 14161 0 net38
rlabel metal2 3450 14756 3450 14756 0 net39
rlabel metal1 1886 11152 1886 11152 0 net4
rlabel metal2 2898 15198 2898 15198 0 net40
rlabel metal2 9982 15572 9982 15572 0 net41
rlabel metal1 1886 17136 1886 17136 0 net42
rlabel metal1 2231 16490 2231 16490 0 net43
rlabel metal1 2346 16762 2346 16762 0 net44
rlabel metal1 14214 8908 14214 8908 0 net45
rlabel metal1 13754 9520 13754 9520 0 net46
rlabel metal1 7498 9656 7498 9656 0 net47
rlabel metal2 12190 9792 12190 9792 0 net48
rlabel metal1 14122 11866 14122 11866 0 net49
rlabel metal1 5336 9146 5336 9146 0 net5
rlabel metal1 13984 12410 13984 12410 0 net50
rlabel metal1 13294 10574 13294 10574 0 net51
rlabel metal1 10856 8602 10856 8602 0 net52
rlabel metal1 14076 15470 14076 15470 0 net53
rlabel via3 9085 2516 9085 2516 0 net54
rlabel metal1 8418 2482 8418 2482 0 net55
rlabel metal1 12972 2958 12972 2958 0 net56
rlabel metal1 12696 5678 12696 5678 0 net57
rlabel metal2 13570 4386 13570 4386 0 net58
rlabel metal2 9890 1700 9890 1700 0 net59
rlabel metal1 2208 8806 2208 8806 0 net6
rlabel metal2 6486 3162 6486 3162 0 net60
rlabel metal1 14076 4182 14076 4182 0 net61
rlabel metal2 13478 3978 13478 3978 0 net62
rlabel metal1 13064 9690 13064 9690 0 net63
rlabel metal1 6440 11186 6440 11186 0 net64
rlabel metal1 1932 5746 1932 5746 0 net65
rlabel metal1 2852 12206 2852 12206 0 net66
rlabel metal1 4968 7378 4968 7378 0 net67
rlabel metal1 8234 13294 8234 13294 0 net68
rlabel metal1 5336 2482 5336 2482 0 net69
rlabel metal1 1242 13906 1242 13906 0 net7
rlabel metal2 8970 4080 8970 4080 0 net70
rlabel metal1 10074 8568 10074 8568 0 net71
rlabel metal1 9752 6222 9752 6222 0 net72
rlabel metal1 12006 7310 12006 7310 0 net73
rlabel metal1 13984 6834 13984 6834 0 net74
rlabel metal2 12742 6528 12742 6528 0 net75
rlabel metal1 6532 2346 6532 2346 0 net76
rlabel metal2 8326 9316 8326 9316 0 net77
rlabel metal1 10150 7786 10150 7786 0 net78
rlabel via1 7677 6698 7677 6698 0 net79
rlabel metal1 1702 1938 1702 1938 0 net8
rlabel metal2 13294 6970 13294 6970 0 net80
rlabel metal1 2238 6698 2238 6698 0 net81
rlabel metal2 5382 12002 5382 12002 0 net82
rlabel metal1 10396 6358 10396 6358 0 net83
rlabel metal1 5653 5678 5653 5678 0 net84
rlabel metal2 7038 3298 7038 3298 0 net85
rlabel metal2 12834 8330 12834 8330 0 net86
rlabel metal2 11454 3944 11454 3944 0 net87
rlabel metal1 8183 8874 8183 8874 0 net88
rlabel metal1 5101 8534 5101 8534 0 net89
rlabel metal1 6624 8942 6624 8942 0 net9
rlabel metal1 10350 6698 10350 6698 0 net90
rlabel metal1 10120 4794 10120 4794 0 net91
rlabel metal1 10483 3094 10483 3094 0 net92
rlabel metal1 11863 8534 11863 8534 0 net93
rlabel metal2 13386 4998 13386 4998 0 net94
rlabel metal1 12052 3162 12052 3162 0 net95
rlabel metal1 13289 6290 13289 6290 0 net96
rlabel metal2 9844 9962 9844 9962 0 net97
rlabel metal1 11316 2550 11316 2550 0 net98
rlabel metal1 9287 13226 9287 13226 0 net99
rlabel metal2 4094 11271 4094 11271 0 prog_clk
rlabel metal1 14674 16558 14674 16558 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 13938 16592 13938 16592 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 16000 20000
<< end >>
