magic
tech sky130A
magscale 1 2
timestamp 1708041250
<< viali >>
rect 9873 9673 9907 9707
rect 10425 9673 10459 9707
rect 2789 9605 2823 9639
rect 2145 9537 2179 9571
rect 2421 9537 2455 9571
rect 9321 9537 9355 9571
rect 9597 9537 9631 9571
rect 10149 9537 10183 9571
rect 9137 9401 9171 9435
rect 1869 9333 1903 9367
rect 1501 9129 1535 9163
rect 9413 9129 9447 9163
rect 9873 9129 9907 9163
rect 10241 9129 10275 9163
rect 2513 9061 2547 9095
rect 2145 8925 2179 8959
rect 2329 8925 2363 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 10057 8925 10091 8959
rect 1777 8857 1811 8891
rect 9597 8857 9631 8891
rect 1961 8789 1995 8823
rect 9137 8789 9171 8823
rect 9413 8585 9447 8619
rect 9873 8585 9907 8619
rect 1777 8449 1811 8483
rect 6009 8449 6043 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 10149 8449 10183 8483
rect 1501 8313 1535 8347
rect 6193 8313 6227 8347
rect 10425 8245 10459 8279
rect 7113 8041 7147 8075
rect 10057 8041 10091 8075
rect 10425 7973 10459 8007
rect 6929 7837 6963 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 9965 7497 9999 7531
rect 1777 7361 1811 7395
rect 9781 7361 9815 7395
rect 9873 7361 9907 7395
rect 10241 7361 10275 7395
rect 1501 7157 1535 7191
rect 9597 7157 9631 7191
rect 10425 7157 10459 7191
rect 8585 6885 8619 6919
rect 9229 6885 9263 6919
rect 9413 6817 9447 6851
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 9597 6749 9631 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 8217 6613 8251 6647
rect 10057 6613 10091 6647
rect 10333 6613 10367 6647
rect 6929 6409 6963 6443
rect 7849 6409 7883 6443
rect 9321 6409 9355 6443
rect 9689 6409 9723 6443
rect 7941 6341 7975 6375
rect 1777 6273 1811 6307
rect 6745 6273 6779 6307
rect 7113 6273 7147 6307
rect 7665 6273 7699 6307
rect 8861 6273 8895 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 10241 6273 10275 6307
rect 8401 6205 8435 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 9965 6137 9999 6171
rect 1501 6069 1535 6103
rect 7297 6069 7331 6103
rect 10425 6069 10459 6103
rect 1961 5865 1995 5899
rect 8677 5865 8711 5899
rect 9137 5865 9171 5899
rect 9781 5729 9815 5763
rect 1777 5661 1811 5695
rect 7113 5661 7147 5695
rect 8585 5661 8619 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 5273 5593 5307 5627
rect 7358 5593 7392 5627
rect 10057 5593 10091 5627
rect 10149 5593 10183 5627
rect 10333 5593 10367 5627
rect 6745 5525 6779 5559
rect 8493 5525 8527 5559
rect 9321 5525 9355 5559
rect 1961 5321 1995 5355
rect 9413 5321 9447 5355
rect 7174 5253 7208 5287
rect 10333 5253 10367 5287
rect 1777 5185 1811 5219
rect 2145 5185 2179 5219
rect 5181 5185 5215 5219
rect 6653 5185 6687 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 9781 5185 9815 5219
rect 5549 5117 5583 5151
rect 6929 5117 6963 5151
rect 8953 5117 8987 5151
rect 9597 5117 9631 5151
rect 10425 5117 10459 5151
rect 6837 5049 6871 5083
rect 8401 5049 8435 5083
rect 1501 4981 1535 5015
rect 5273 4981 5307 5015
rect 6193 4981 6227 5015
rect 8309 4981 8343 5015
rect 1777 4777 1811 4811
rect 4353 4777 4387 4811
rect 7113 4777 7147 4811
rect 5733 4641 5767 4675
rect 8309 4641 8343 4675
rect 1593 4573 1627 4607
rect 5477 4573 5511 4607
rect 7665 4573 7699 4607
rect 8401 4573 8435 4607
rect 9689 4573 9723 4607
rect 10057 4573 10091 4607
rect 10149 4573 10183 4607
rect 5825 4505 5859 4539
rect 8585 4437 8619 4471
rect 9137 4437 9171 4471
rect 9873 4437 9907 4471
rect 10241 4437 10275 4471
rect 2329 4233 2363 4267
rect 4997 4233 5031 4267
rect 8677 4233 8711 4267
rect 9597 4233 9631 4267
rect 5641 4165 5675 4199
rect 7564 4165 7598 4199
rect 1777 4097 1811 4131
rect 2237 4097 2271 4131
rect 2513 4097 2547 4131
rect 2605 4097 2639 4131
rect 3709 4097 3743 4131
rect 4813 4097 4847 4131
rect 7297 4097 7331 4131
rect 9689 4097 9723 4131
rect 3985 4029 4019 4063
rect 5457 4029 5491 4063
rect 5733 4029 5767 4063
rect 5917 4029 5951 4063
rect 7113 4029 7147 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 9873 4029 9907 4063
rect 3893 3961 3927 3995
rect 1501 3893 1535 3927
rect 2053 3893 2087 3927
rect 2789 3893 2823 3927
rect 4629 3893 4663 3927
rect 6561 3893 6595 3927
rect 10241 3893 10275 3927
rect 1961 3689 1995 3723
rect 2421 3689 2455 3723
rect 2697 3689 2731 3723
rect 3617 3689 3651 3723
rect 5457 3689 5491 3723
rect 6929 3689 6963 3723
rect 9965 3621 9999 3655
rect 5917 3553 5951 3587
rect 1409 3485 1443 3519
rect 2053 3485 2087 3519
rect 2329 3485 2363 3519
rect 2605 3485 2639 3519
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 6377 3485 6411 3519
rect 6837 3485 6871 3519
rect 8042 3485 8076 3519
rect 8309 3485 8343 3519
rect 8769 3485 8803 3519
rect 9505 3485 9539 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 4344 3417 4378 3451
rect 5641 3417 5675 3451
rect 5733 3417 5767 3451
rect 1593 3349 1627 3383
rect 2237 3349 2271 3383
rect 3249 3349 3283 3383
rect 3893 3349 3927 3383
rect 6469 3349 6503 3383
rect 6653 3349 6687 3383
rect 8585 3349 8619 3383
rect 8953 3349 8987 3383
rect 1961 3145 1995 3179
rect 2421 3145 2455 3179
rect 3249 3145 3283 3179
rect 3617 3145 3651 3179
rect 7297 3145 7331 3179
rect 9045 3145 9079 3179
rect 10425 3145 10459 3179
rect 1777 3077 1811 3111
rect 4752 3077 4786 3111
rect 6561 3077 6595 3111
rect 7113 3077 7147 3111
rect 7748 3077 7782 3111
rect 10057 3077 10091 3111
rect 10149 3077 10183 3111
rect 2145 3009 2179 3043
rect 2237 3009 2271 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 8953 3009 8987 3043
rect 9413 3009 9447 3043
rect 10333 3009 10367 3043
rect 4997 2941 5031 2975
rect 6193 2941 6227 2975
rect 6469 2941 6503 2975
rect 2697 2873 2731 2907
rect 3341 2873 3375 2907
rect 9597 2873 9631 2907
rect 1501 2805 1535 2839
rect 2973 2805 3007 2839
rect 5365 2805 5399 2839
rect 8861 2805 8895 2839
rect 9229 2805 9263 2839
rect 2697 2601 2731 2635
rect 4169 2601 4203 2635
rect 4905 2601 4939 2635
rect 7021 2601 7055 2635
rect 7389 2601 7423 2635
rect 8677 2601 8711 2635
rect 9597 2601 9631 2635
rect 10333 2601 10367 2635
rect 1869 2533 1903 2567
rect 6653 2533 6687 2567
rect 2053 2465 2087 2499
rect 2973 2465 3007 2499
rect 3157 2465 3191 2499
rect 3617 2465 3651 2499
rect 8401 2465 8435 2499
rect 9689 2465 9723 2499
rect 9873 2465 9907 2499
rect 1593 2397 1627 2431
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 2881 2397 2915 2431
rect 3893 2397 3927 2431
rect 4353 2397 4387 2431
rect 6193 2397 6227 2431
rect 6469 2397 6503 2431
rect 6837 2397 6871 2431
rect 7297 2397 7331 2431
rect 7573 2397 7607 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 8953 2397 8987 2431
rect 9137 2397 9171 2431
rect 1501 2261 1535 2295
rect 2605 2261 2639 2295
rect 4077 2261 4111 2295
rect 7113 2261 7147 2295
rect 7757 2261 7791 2295
rect 8033 2261 8067 2295
<< metal1 >>
rect 1104 9818 11016 9840
rect 1104 9766 3388 9818
rect 3440 9766 3452 9818
rect 3504 9766 3516 9818
rect 3568 9766 3580 9818
rect 3632 9766 3644 9818
rect 3696 9766 5826 9818
rect 5878 9766 5890 9818
rect 5942 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 8264 9818
rect 8316 9766 8328 9818
rect 8380 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 10702 9818
rect 10754 9766 10766 9818
rect 10818 9766 10830 9818
rect 10882 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11016 9818
rect 1104 9744 11016 9766
rect 9861 9707 9919 9713
rect 9861 9673 9873 9707
rect 9907 9704 9919 9707
rect 9950 9704 9956 9716
rect 9907 9676 9956 9704
rect 9907 9673 9919 9676
rect 9861 9667 9919 9673
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10413 9707 10471 9713
rect 10413 9673 10425 9707
rect 10459 9704 10471 9707
rect 10502 9704 10508 9716
rect 10459 9676 10508 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 2774 9596 2780 9648
rect 2832 9596 2838 9648
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1912 9540 2145 9568
rect 1912 9528 1918 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2424 9500 2452 9531
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9456 9540 9597 9568
rect 9456 9528 9462 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 2004 9472 2452 9500
rect 2004 9460 2010 9472
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9214 9432 9220 9444
rect 9171 9404 9220 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 992 9336 1869 9364
rect 992 9324 998 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 1486 9120 1492 9172
rect 1544 9120 1550 9172
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 10042 9160 10048 9172
rect 9907 9132 10048 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10226 9120 10232 9172
rect 10284 9120 10290 9172
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 10134 9092 10140 9104
rect 2547 9064 10140 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8888 1823 8891
rect 2148 8888 2176 8919
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 4304 8928 8953 8956
rect 4304 8916 4310 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8941 8919 8999 8925
rect 9048 8928 9229 8956
rect 4522 8888 4528 8900
rect 1811 8860 1992 8888
rect 2148 8860 4528 8888
rect 1811 8857 1823 8860
rect 1765 8851 1823 8857
rect 1964 8829 1992 8860
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8789 2007 8823
rect 1949 8783 2007 8789
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 9048 8820 9076 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 9140 8860 9597 8888
rect 9140 8829 9168 8860
rect 9585 8857 9597 8860
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 2924 8792 9076 8820
rect 9125 8823 9183 8829
rect 2924 8780 2930 8792
rect 9125 8789 9137 8823
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 1104 8730 11016 8752
rect 1104 8678 3388 8730
rect 3440 8678 3452 8730
rect 3504 8678 3516 8730
rect 3568 8678 3580 8730
rect 3632 8678 3644 8730
rect 3696 8678 5826 8730
rect 5878 8678 5890 8730
rect 5942 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 8264 8730
rect 8316 8678 8328 8730
rect 8380 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 10702 8730
rect 10754 8678 10766 8730
rect 10818 8678 10830 8730
rect 10882 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11016 8730
rect 1104 8656 11016 8678
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 9364 8588 9413 8616
rect 9364 8576 9370 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 9861 8619 9919 8625
rect 9861 8585 9873 8619
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 9876 8548 9904 8579
rect 10594 8548 10600 8560
rect 9876 8520 10600 8548
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2038 8480 2044 8492
rect 1811 8452 2044 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 3936 8452 6009 8480
rect 3936 8440 3942 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 5997 8443 6055 8449
rect 6886 8452 9597 8480
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 6886 8412 6914 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 2832 8384 6914 8412
rect 2832 8372 2838 8384
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 9692 8344 9720 8443
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9916 8452 10149 8480
rect 9916 8440 9922 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 6227 8316 9720 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 10502 8276 10508 8288
rect 10459 8248 10508 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 9858 8072 9864 8084
rect 7147 8044 9864 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10042 8032 10048 8084
rect 10100 8032 10106 8084
rect 10410 7964 10416 8016
rect 10468 7964 10474 8016
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7466 7868 7472 7880
rect 6963 7840 7472 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 8996 7840 9873 7868
rect 8996 7828 9002 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 1104 7642 11016 7664
rect 1104 7590 3388 7642
rect 3440 7590 3452 7642
rect 3504 7590 3516 7642
rect 3568 7590 3580 7642
rect 3632 7590 3644 7642
rect 3696 7590 5826 7642
rect 5878 7590 5890 7642
rect 5942 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 8264 7642
rect 8316 7590 8328 7642
rect 8380 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 10702 7642
rect 10754 7590 10766 7642
rect 10818 7590 10830 7642
rect 10882 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11016 7642
rect 1104 7568 11016 7590
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10226 7528 10232 7540
rect 9999 7500 10232 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 9364 7432 9904 7460
rect 9364 7420 9370 7432
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2590 7392 2596 7404
rect 1811 7364 2596 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 9876 7401 9904 7432
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9784 7324 9812 7355
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 10502 7324 10508 7336
rect 9784 7296 10508 7324
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 6880 7160 9597 7188
rect 6880 7148 6886 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 10410 7148 10416 7200
rect 10468 7148 10474 7200
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 8588 6956 9444 6984
rect 8588 6925 8616 6956
rect 8573 6919 8631 6925
rect 8573 6885 8585 6919
rect 8619 6885 8631 6919
rect 8573 6879 8631 6885
rect 9217 6919 9275 6925
rect 9217 6885 9229 6919
rect 9263 6916 9275 6919
rect 9306 6916 9312 6928
rect 9263 6888 9312 6916
rect 9263 6885 9275 6888
rect 9217 6879 9275 6885
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 9416 6857 9444 6956
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9631 6752 9689 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 8404 6712 8432 6743
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10008 6752 10241 6780
rect 10008 6740 10014 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10870 6780 10876 6792
rect 10551 6752 10876 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 7892 6684 8432 6712
rect 7892 6672 7898 6684
rect 8205 6647 8263 6653
rect 8205 6613 8217 6647
rect 8251 6644 8263 6647
rect 8754 6644 8760 6656
rect 8251 6616 8760 6644
rect 8251 6613 8263 6616
rect 8205 6607 8263 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 10042 6604 10048 6656
rect 10100 6604 10106 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10192 6616 10333 6644
rect 10192 6604 10198 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 1104 6554 11016 6576
rect 1104 6502 3388 6554
rect 3440 6502 3452 6554
rect 3504 6502 3516 6554
rect 3568 6502 3580 6554
rect 3632 6502 3644 6554
rect 3696 6502 5826 6554
rect 5878 6502 5890 6554
rect 5942 6502 5954 6554
rect 6006 6502 6018 6554
rect 6070 6502 6082 6554
rect 6134 6502 8264 6554
rect 8316 6502 8328 6554
rect 8380 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 10702 6554
rect 10754 6502 10766 6554
rect 10818 6502 10830 6554
rect 10882 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11016 6554
rect 1104 6480 11016 6502
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6409 6975 6443
rect 6917 6403 6975 6409
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6730 6304 6736 6316
rect 5592 6276 6736 6304
rect 5592 6264 5598 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 6932 6304 6960 6403
rect 7834 6400 7840 6452
rect 7892 6400 7898 6452
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 10226 6440 10232 6452
rect 9723 6412 10232 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6372 7987 6375
rect 7975 6344 8708 6372
rect 7975 6341 7987 6344
rect 7929 6335 7987 6341
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6932 6276 7113 6304
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 8110 6304 8116 6316
rect 7699 6276 8116 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 8110 6264 8116 6276
rect 8168 6304 8174 6316
rect 8168 6276 8524 6304
rect 8168 6264 8174 6276
rect 8496 6248 8524 6276
rect 8386 6196 8392 6248
rect 8444 6196 8450 6248
rect 8478 6196 8484 6248
rect 8536 6196 8542 6248
rect 8680 6245 8708 6344
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9088 6344 10272 6372
rect 9088 6332 9094 6344
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8812 6276 8861 6304
rect 8812 6264 8818 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 10134 6304 10140 6316
rect 10091 6276 10140 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10244 6313 10272 6344
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9214 6236 9220 6248
rect 8711 6208 9220 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 8588 6168 8616 6199
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 8588 6140 9965 6168
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 934 6060 940 6112
rect 992 6100 998 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 992 6072 1501 6100
rect 992 6060 998 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1489 6063 1547 6069
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7834 6100 7840 6112
rect 7331 6072 7840 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 1946 5856 1952 5908
rect 2004 5856 2010 5908
rect 6822 5896 6828 5908
rect 2746 5868 6828 5896
rect 2746 5828 2774 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8444 5868 8677 5896
rect 8444 5856 8450 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9950 5896 9956 5908
rect 9171 5868 9956 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 1780 5800 2774 5828
rect 1780 5701 1808 5800
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 6788 5732 7236 5760
rect 6788 5720 6794 5732
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 1765 5655 1823 5661
rect 6932 5664 7113 5692
rect 5261 5627 5319 5633
rect 5261 5593 5273 5627
rect 5307 5624 5319 5627
rect 6178 5624 6184 5636
rect 5307 5596 6184 5624
rect 5307 5593 5319 5596
rect 5261 5587 5319 5593
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 6932 5568 6960 5664
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 7208 5692 7236 5732
rect 9766 5720 9772 5772
rect 9824 5720 9830 5772
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 7208 5664 8585 5692
rect 7101 5655 7159 5661
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8812 5664 8953 5692
rect 8812 5652 8818 5664
rect 8941 5661 8953 5664
rect 8987 5692 8999 5695
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8987 5664 9229 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 7346 5627 7404 5633
rect 7346 5624 7358 5627
rect 7248 5596 7358 5624
rect 7248 5584 7254 5596
rect 7346 5593 7358 5596
rect 7392 5593 7404 5627
rect 7346 5587 7404 5593
rect 10042 5584 10048 5636
rect 10100 5584 10106 5636
rect 10137 5627 10195 5633
rect 10137 5593 10149 5627
rect 10183 5624 10195 5627
rect 10321 5627 10379 5633
rect 10321 5624 10333 5627
rect 10183 5596 10333 5624
rect 10183 5593 10195 5596
rect 10137 5587 10195 5593
rect 10321 5593 10333 5596
rect 10367 5593 10379 5627
rect 10321 5587 10379 5593
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5556 6791 5559
rect 6914 5556 6920 5568
rect 6779 5528 6920 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8938 5556 8944 5568
rect 8536 5528 8944 5556
rect 8536 5516 8542 5528
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 1104 5466 11016 5488
rect 1104 5414 3388 5466
rect 3440 5414 3452 5466
rect 3504 5414 3516 5466
rect 3568 5414 3580 5466
rect 3632 5414 3644 5466
rect 3696 5414 5826 5466
rect 5878 5414 5890 5466
rect 5942 5414 5954 5466
rect 6006 5414 6018 5466
rect 6070 5414 6082 5466
rect 6134 5414 8264 5466
rect 8316 5414 8328 5466
rect 8380 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 10702 5466
rect 10754 5414 10766 5466
rect 10818 5414 10830 5466
rect 10882 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11016 5466
rect 1104 5392 11016 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1820 5324 1961 5352
rect 1820 5312 1826 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 5442 5352 5448 5364
rect 1949 5315 2007 5321
rect 5184 5324 5448 5352
rect 1762 5176 1768 5228
rect 1820 5176 1826 5228
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 1872 5188 2145 5216
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 1872 5148 1900 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 5184 5225 5212 5324
rect 5442 5312 5448 5324
rect 5500 5352 5506 5364
rect 9030 5352 9036 5364
rect 5500 5324 9036 5352
rect 5500 5312 5506 5324
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 10410 5352 10416 5364
rect 9447 5324 10416 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 6822 5244 6828 5296
rect 6880 5284 6886 5296
rect 7162 5287 7220 5293
rect 7162 5284 7174 5287
rect 6880 5256 7174 5284
rect 6880 5244 6886 5256
rect 7162 5253 7174 5256
rect 7208 5253 7220 5287
rect 7162 5247 7220 5253
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 10321 5287 10379 5293
rect 10321 5284 10333 5287
rect 9364 5256 10333 5284
rect 9364 5244 9370 5256
rect 10321 5253 10333 5256
rect 10367 5253 10379 5287
rect 10321 5247 10379 5253
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4212 5188 5181 5216
rect 4212 5176 4218 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 9030 5216 9036 5228
rect 6687 5188 9036 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 9217 5179 9275 5185
rect 9324 5188 9505 5216
rect 1728 5120 1900 5148
rect 1728 5108 1734 5120
rect 4338 5108 4344 5160
rect 4396 5148 4402 5160
rect 5534 5148 5540 5160
rect 4396 5120 5540 5148
rect 4396 5108 4402 5120
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 6914 5108 6920 5160
rect 6972 5108 6978 5160
rect 8938 5108 8944 5160
rect 8996 5108 9002 5160
rect 6822 5040 6828 5092
rect 6880 5040 6886 5092
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 8168 5052 8401 5080
rect 8168 5040 8174 5052
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 9232 5080 9260 5179
rect 9324 5160 9352 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 9306 5108 9312 5160
rect 9364 5108 9370 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 9456 5120 9597 5148
rect 9456 5108 9462 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 9585 5111 9643 5117
rect 10336 5120 10425 5148
rect 10226 5080 10232 5092
rect 9232 5052 10232 5080
rect 8389 5043 8447 5049
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10336 5024 10364 5120
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 5261 5015 5319 5021
rect 5261 4981 5273 5015
rect 5307 5012 5319 5015
rect 5718 5012 5724 5024
rect 5307 4984 5724 5012
rect 5307 4981 5319 4984
rect 5261 4975 5319 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 7190 5012 7196 5024
rect 6227 4984 7196 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 8294 4972 8300 5024
rect 8352 4972 8358 5024
rect 10318 4972 10324 5024
rect 10376 4972 10382 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 4246 4808 4252 4820
rect 1811 4780 4252 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 4338 4768 4344 4820
rect 4396 4768 4402 4820
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 7101 4811 7159 4817
rect 7101 4808 7113 4811
rect 6236 4780 7113 4808
rect 6236 4768 6242 4780
rect 7101 4777 7113 4780
rect 7147 4777 7159 4811
rect 7101 4771 7159 4777
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7064 4712 10180 4740
rect 7064 4700 7070 4712
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6914 4672 6920 4684
rect 5767 4644 6920 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6914 4632 6920 4644
rect 6972 4672 6978 4684
rect 7282 4672 7288 4684
rect 6972 4644 7288 4672
rect 6972 4632 6978 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8754 4672 8760 4684
rect 8343 4644 8760 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 1946 4604 1952 4616
rect 1627 4576 1952 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 5465 4607 5523 4613
rect 5465 4573 5477 4607
rect 5511 4604 5523 4607
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 5511 4576 7665 4604
rect 5511 4573 5523 4576
rect 5465 4567 5523 4573
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 7653 4567 7711 4573
rect 8312 4576 8401 4604
rect 8312 4548 8340 4576
rect 8389 4573 8401 4576
rect 8435 4604 8447 4607
rect 9030 4604 9036 4616
rect 8435 4576 9036 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 9030 4564 9036 4576
rect 9088 4604 9094 4616
rect 10152 4613 10180 4712
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9088 4576 9689 4604
rect 9088 4564 9094 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 5813 4539 5871 4545
rect 5813 4505 5825 4539
rect 5859 4505 5871 4539
rect 5813 4499 5871 4505
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 5828 4468 5856 4499
rect 8294 4496 8300 4548
rect 8352 4496 8358 4548
rect 10060 4536 10088 4567
rect 8588 4508 10088 4536
rect 8588 4477 8616 4508
rect 4488 4440 5856 4468
rect 8573 4471 8631 4477
rect 4488 4428 4494 4440
rect 8573 4437 8585 4471
rect 8619 4437 8631 4471
rect 8573 4431 8631 4437
rect 9122 4428 9128 4480
rect 9180 4428 9186 4480
rect 9858 4428 9864 4480
rect 9916 4428 9922 4480
rect 10226 4428 10232 4480
rect 10284 4428 10290 4480
rect 1104 4378 11016 4400
rect 1104 4326 3388 4378
rect 3440 4326 3452 4378
rect 3504 4326 3516 4378
rect 3568 4326 3580 4378
rect 3632 4326 3644 4378
rect 3696 4326 5826 4378
rect 5878 4326 5890 4378
rect 5942 4326 5954 4378
rect 6006 4326 6018 4378
rect 6070 4326 6082 4378
rect 6134 4326 8264 4378
rect 8316 4326 8328 4378
rect 8380 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 10702 4378
rect 10754 4326 10766 4378
rect 10818 4326 10830 4378
rect 10882 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11016 4378
rect 1104 4304 11016 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 2317 4267 2375 4273
rect 2317 4264 2329 4267
rect 1820 4236 2329 4264
rect 1820 4224 1826 4236
rect 2317 4233 2329 4236
rect 2363 4233 2375 4267
rect 2317 4227 2375 4233
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4948 4236 4997 4264
rect 4948 4224 4954 4236
rect 4985 4233 4997 4236
rect 5031 4233 5043 4267
rect 4985 4227 5043 4233
rect 8665 4267 8723 4273
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 8754 4264 8760 4276
rect 8711 4236 8760 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9272 4236 9597 4264
rect 9272 4224 9278 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 4154 4196 4160 4208
rect 3712 4168 4160 4196
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 2222 4088 2228 4140
rect 2280 4088 2286 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 3142 4128 3148 4140
rect 2639 4100 3148 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2516 4060 2544 4091
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3712 4137 3740 4168
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 5258 4156 5264 4208
rect 5316 4196 5322 4208
rect 5629 4199 5687 4205
rect 5629 4196 5641 4199
rect 5316 4168 5641 4196
rect 5316 4156 5322 4168
rect 5629 4165 5641 4168
rect 5675 4165 5687 4199
rect 5629 4159 5687 4165
rect 7552 4199 7610 4205
rect 7552 4165 7564 4199
rect 7598 4196 7610 4199
rect 9122 4196 9128 4208
rect 7598 4168 9128 4196
rect 7598 4165 7610 4168
rect 7552 4159 7610 4165
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 3697 4091 3755 4097
rect 3896 4100 4813 4128
rect 2682 4060 2688 4072
rect 2516 4032 2688 4060
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3896 4001 3924 4100
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 9677 4131 9735 4137
rect 7892 4100 9168 4128
rect 7892 4088 7898 4100
rect 3970 4020 3976 4072
rect 4028 4020 4034 4072
rect 5350 4060 5356 4072
rect 4080 4032 5356 4060
rect 3881 3995 3939 4001
rect 3881 3961 3893 3995
rect 3927 3961 3939 3995
rect 4080 3992 4108 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5721 4063 5779 4069
rect 5491 4032 5672 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5644 4004 5672 4032
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5767 4032 5917 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 7098 4060 7104 4072
rect 6604 4032 7104 4060
rect 6604 4020 6610 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9140 4069 9168 4100
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 10226 4128 10232 4140
rect 9723 4100 10232 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8720 4032 8953 4060
rect 8720 4020 8726 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9364 4032 9873 4060
rect 9364 4020 9370 4032
rect 9861 4029 9873 4032
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 5626 3992 5632 4004
rect 3881 3955 3939 3961
rect 3988 3964 4108 3992
rect 4356 3964 5632 3992
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 992 3896 1501 3924
rect 992 3884 998 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 2038 3884 2044 3936
rect 2096 3884 2102 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 3988 3924 4016 3964
rect 3016 3896 4016 3924
rect 3016 3884 3022 3896
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4356 3924 4384 3964
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 4120 3896 4384 3924
rect 4120 3884 4126 3896
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4488 3896 4629 3924
rect 4488 3884 4494 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5408 3896 6561 3924
rect 5408 3884 5414 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 8846 3924 8852 3936
rect 6788 3896 8852 3924
rect 6788 3884 6794 3896
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 10226 3884 10232 3936
rect 10284 3884 10290 3936
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1820 3692 1961 3720
rect 1820 3680 1826 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2498 3720 2504 3732
rect 2455 3692 2504 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2648 3692 2697 3720
rect 2648 3680 2654 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3878 3720 3884 3732
rect 3651 3692 3884 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5442 3680 5448 3732
rect 5500 3680 5506 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6730 3720 6736 3732
rect 5592 3692 6736 3720
rect 5592 3680 5598 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 6917 3723 6975 3729
rect 6917 3689 6929 3723
rect 6963 3720 6975 3723
rect 7006 3720 7012 3732
rect 6963 3692 7012 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 7006 3680 7012 3692
rect 7064 3720 7070 3732
rect 7064 3692 8892 3720
rect 7064 3680 7070 3692
rect 4062 3652 4068 3664
rect 2056 3624 4068 3652
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 2056 3525 2084 3624
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 3970 3584 3976 3596
rect 2746 3556 3976 3584
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 900 3488 1409 3516
rect 900 3476 906 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2314 3476 2320 3528
rect 2372 3476 2378 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2608 3448 2636 3479
rect 2004 3420 2636 3448
rect 2004 3408 2010 3420
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 1762 3380 1768 3392
rect 1627 3352 1768 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 2406 3340 2412 3392
rect 2464 3380 2470 3392
rect 2746 3380 2774 3556
rect 3804 3528 3832 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5684 3556 5917 3584
rect 5684 3544 5690 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 8864 3528 8892 3692
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3652 10011 3655
rect 10134 3652 10140 3664
rect 9999 3624 10140 3652
rect 9999 3621 10011 3624
rect 9953 3615 10011 3621
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 2866 3476 2872 3528
rect 2924 3476 2930 3528
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3436 3448 3464 3479
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 6365 3519 6423 3525
rect 4111 3488 5028 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4332 3451 4390 3457
rect 3436 3420 4154 3448
rect 2464 3352 2774 3380
rect 2464 3340 2470 3352
rect 3234 3340 3240 3392
rect 3292 3340 3298 3392
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 4126 3380 4154 3420
rect 4332 3417 4344 3451
rect 4378 3448 4390 3451
rect 4430 3448 4436 3460
rect 4378 3420 4436 3448
rect 4378 3417 4390 3420
rect 4332 3411 4390 3417
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 5000 3392 5028 3488
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 5626 3408 5632 3460
rect 5684 3408 5690 3460
rect 5718 3408 5724 3460
rect 5776 3408 5782 3460
rect 4614 3380 4620 3392
rect 4126 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4982 3340 4988 3392
rect 5040 3340 5046 3392
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 6380 3380 6408 3479
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 8030 3519 8088 3525
rect 8030 3485 8042 3519
rect 8076 3485 8088 3519
rect 8030 3479 8088 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8036 3448 8064 3479
rect 8110 3448 8116 3460
rect 8036 3420 8116 3448
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 5316 3352 6408 3380
rect 5316 3340 5322 3352
rect 6454 3340 6460 3392
rect 6512 3340 6518 3392
rect 6638 3340 6644 3392
rect 6696 3340 6702 3392
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 8312 3380 8340 3479
rect 8772 3448 8800 3479
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 8904 3488 9505 3516
rect 8904 3476 8910 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9640 3488 10149 3516
rect 9640 3476 9646 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10318 3476 10324 3528
rect 10376 3476 10382 3528
rect 11054 3448 11060 3460
rect 8772 3420 11060 3448
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 7616 3352 8340 3380
rect 7616 3340 7622 3352
rect 8570 3340 8576 3392
rect 8628 3340 8634 3392
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 1104 3290 11016 3312
rect 1104 3238 3388 3290
rect 3440 3238 3452 3290
rect 3504 3238 3516 3290
rect 3568 3238 3580 3290
rect 3632 3238 3644 3290
rect 3696 3238 5826 3290
rect 5878 3238 5890 3290
rect 5942 3238 5954 3290
rect 6006 3238 6018 3290
rect 6070 3238 6082 3290
rect 6134 3238 8264 3290
rect 8316 3238 8328 3290
rect 8380 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 10702 3290
rect 10754 3238 10766 3290
rect 10818 3238 10830 3290
rect 10882 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11016 3290
rect 1104 3216 11016 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1912 3148 1961 3176
rect 1912 3136 1918 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 3050 3176 3056 3188
rect 2455 3148 3056 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3326 3176 3332 3188
rect 3283 3148 3332 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 3786 3176 3792 3188
rect 3651 3148 3792 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 3936 3148 5580 3176
rect 3936 3136 3942 3148
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 2240 3108 2268 3136
rect 4522 3108 4528 3120
rect 1811 3080 2268 3108
rect 2516 3080 4528 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 2130 3000 2136 3052
rect 2188 3000 2194 3052
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2406 3040 2412 3052
rect 2271 3012 2412 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2516 3049 2544 3080
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4614 3068 4620 3120
rect 4672 3068 4678 3120
rect 4740 3111 4798 3117
rect 4740 3077 4752 3111
rect 4786 3108 4798 3111
rect 5350 3108 5356 3120
rect 4786 3080 5356 3108
rect 4786 3077 4798 3080
rect 4740 3071 4798 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 2958 3040 2964 3052
rect 2823 3012 2964 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3513 3043 3571 3049
rect 3099 3012 3372 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3344 2913 3372 3012
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 4430 3040 4436 3052
rect 3559 3012 4436 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4632 3040 4660 3068
rect 5442 3040 5448 3052
rect 4632 3012 5448 3040
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5552 3049 5580 3148
rect 6454 3136 6460 3188
rect 6512 3136 6518 3188
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 8662 3176 8668 3188
rect 7331 3148 8668 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 8938 3136 8944 3188
rect 8996 3136 9002 3188
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9306 3176 9312 3188
rect 9079 3148 9312 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9456 3148 10088 3176
rect 9456 3136 9462 3148
rect 6472 3108 6500 3136
rect 5736 3080 6500 3108
rect 6549 3111 6607 3117
rect 5736 3049 5764 3080
rect 6549 3077 6561 3111
rect 6595 3108 6607 3111
rect 6638 3108 6644 3120
rect 6595 3080 6644 3108
rect 6595 3077 6607 3080
rect 6549 3071 6607 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 6788 3080 7113 3108
rect 6788 3068 6794 3080
rect 7101 3077 7113 3080
rect 7147 3108 7159 3111
rect 7736 3111 7794 3117
rect 7147 3080 7696 3108
rect 7147 3077 7159 3080
rect 7101 3071 7159 3077
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7558 3040 7564 3052
rect 7515 3012 7564 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6457 2975 6515 2981
rect 6457 2972 6469 2975
rect 6227 2944 6469 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6457 2941 6469 2944
rect 6503 2941 6515 2975
rect 7484 2972 7512 3003
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 7668 3040 7696 3080
rect 7736 3077 7748 3111
rect 7782 3108 7794 3111
rect 8956 3108 8984 3136
rect 10060 3117 10088 3148
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10376 3148 10425 3176
rect 10376 3136 10382 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 7782 3080 8984 3108
rect 10045 3111 10103 3117
rect 7782 3077 7794 3080
rect 7736 3071 7794 3077
rect 10045 3077 10057 3111
rect 10091 3077 10103 3111
rect 10045 3071 10103 3077
rect 10134 3068 10140 3120
rect 10192 3068 10198 3120
rect 8941 3043 8999 3049
rect 7668 3012 8524 3040
rect 6457 2935 6515 2941
rect 6886 2944 7512 2972
rect 8496 2972 8524 3012
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9030 3040 9036 3052
rect 8987 3012 9036 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 10410 3040 10416 3052
rect 10367 3012 10416 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 9416 2972 9444 3003
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10502 2972 10508 2984
rect 8496 2944 9352 2972
rect 9416 2944 10508 2972
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2648 2876 2697 2904
rect 2648 2864 2654 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 2685 2867 2743 2873
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2873 3387 2907
rect 3329 2867 3387 2873
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 6886 2904 6914 2944
rect 9324 2904 9352 2944
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 9585 2907 9643 2913
rect 9585 2904 9597 2907
rect 5132 2876 6914 2904
rect 7208 2876 7420 2904
rect 5132 2864 5138 2876
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 5258 2836 5264 2848
rect 3007 2808 5264 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5353 2839 5411 2845
rect 5353 2805 5365 2839
rect 5399 2836 5411 2839
rect 5626 2836 5632 2848
rect 5399 2808 5632 2836
rect 5399 2805 5411 2808
rect 5353 2799 5411 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 7208 2836 7236 2876
rect 6328 2808 7236 2836
rect 7392 2836 7420 2876
rect 8404 2876 9260 2904
rect 9324 2876 9597 2904
rect 8404 2836 8432 2876
rect 7392 2808 8432 2836
rect 8849 2839 8907 2845
rect 6328 2796 6334 2808
rect 8849 2805 8861 2839
rect 8895 2836 8907 2839
rect 9122 2836 9128 2848
rect 8895 2808 9128 2836
rect 8895 2805 8907 2808
rect 8849 2799 8907 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9232 2845 9260 2876
rect 9585 2873 9597 2876
rect 9631 2873 9643 2907
rect 9585 2867 9643 2873
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2805 9275 2839
rect 9217 2799 9275 2805
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 2682 2592 2688 2644
rect 2740 2592 2746 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4338 2632 4344 2644
rect 4203 2604 4344 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5074 2632 5080 2644
rect 4939 2604 5080 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 6822 2632 6828 2644
rect 5491 2604 6828 2632
rect 1857 2567 1915 2573
rect 1857 2533 1869 2567
rect 1903 2564 1915 2567
rect 5491 2564 5519 2604
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7009 2635 7067 2641
rect 7009 2632 7021 2635
rect 6972 2604 7021 2632
rect 6972 2592 6978 2604
rect 7009 2601 7021 2604
rect 7055 2601 7067 2635
rect 7009 2595 7067 2601
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9398 2632 9404 2644
rect 8711 2604 9404 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9585 2635 9643 2641
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10134 2632 10140 2644
rect 9631 2604 10140 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10318 2592 10324 2644
rect 10376 2592 10382 2644
rect 1903 2536 5519 2564
rect 6641 2567 6699 2573
rect 1903 2533 1915 2536
rect 1857 2527 1915 2533
rect 6641 2533 6653 2567
rect 6687 2564 6699 2567
rect 7466 2564 7472 2576
rect 6687 2536 7472 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 2961 2499 3019 2505
rect 2961 2496 2973 2499
rect 2087 2468 2973 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 2961 2465 2973 2468
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 3142 2456 3148 2508
rect 3200 2456 3206 2508
rect 3605 2499 3663 2505
rect 3605 2465 3617 2499
rect 3651 2496 3663 2499
rect 5626 2496 5632 2508
rect 3651 2468 5632 2496
rect 3651 2465 3663 2468
rect 3605 2459 3663 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 7006 2496 7012 2508
rect 6104 2468 7012 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1596 2360 1624 2391
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1820 2400 1961 2428
rect 1820 2388 1826 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2406 2388 2412 2440
rect 2464 2388 2470 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3786 2428 3792 2440
rect 2915 2400 3792 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 6104 2428 6132 2468
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 8389 2499 8447 2505
rect 7300 2468 8156 2496
rect 4387 2400 6132 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 6454 2388 6460 2440
rect 6512 2388 6518 2440
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 6914 2428 6920 2440
rect 6871 2400 6920 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7300 2437 7328 2468
rect 8128 2440 8156 2468
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 8435 2468 9689 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 9858 2456 9864 2508
rect 9916 2456 9922 2508
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 7944 2360 7972 2391
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8846 2428 8852 2440
rect 8619 2400 8852 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 10042 2360 10048 2372
rect 1596 2332 7788 2360
rect 7944 2332 10048 2360
rect 1486 2252 1492 2304
rect 1544 2252 1550 2304
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2292 2651 2295
rect 2774 2292 2780 2304
rect 2639 2264 2780 2292
rect 2639 2261 2651 2264
rect 2593 2255 2651 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 4065 2295 4123 2301
rect 4065 2261 4077 2295
rect 4111 2292 4123 2295
rect 5534 2292 5540 2304
rect 4111 2264 5540 2292
rect 4111 2261 4123 2264
rect 4065 2255 4123 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 7760 2301 7788 2332
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2261 7803 2295
rect 7745 2255 7803 2261
rect 8018 2252 8024 2304
rect 8076 2252 8082 2304
rect 1104 2202 11016 2224
rect 1104 2150 3388 2202
rect 3440 2150 3452 2202
rect 3504 2150 3516 2202
rect 3568 2150 3580 2202
rect 3632 2150 3644 2202
rect 3696 2150 5826 2202
rect 5878 2150 5890 2202
rect 5942 2150 5954 2202
rect 6006 2150 6018 2202
rect 6070 2150 6082 2202
rect 6134 2150 8264 2202
rect 8316 2150 8328 2202
rect 8380 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 10702 2202
rect 10754 2150 10766 2202
rect 10818 2150 10830 2202
rect 10882 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11016 2202
rect 1104 2128 11016 2150
rect 1486 2048 1492 2100
rect 1544 2048 1550 2100
rect 2958 2048 2964 2100
rect 3016 2088 3022 2100
rect 7098 2088 7104 2100
rect 3016 2060 7104 2088
rect 3016 2048 3022 2060
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 1504 1952 1532 2048
rect 3878 1980 3884 2032
rect 3936 2020 3942 2032
rect 8202 2020 8208 2032
rect 3936 1992 8208 2020
rect 3936 1980 3942 1992
rect 8202 1980 8208 1992
rect 8260 1980 8266 2032
rect 1504 1924 2774 1952
rect 1670 1844 1676 1896
rect 1728 1844 1734 1896
rect 2746 1884 2774 1924
rect 2746 1856 3004 1884
rect 1688 1816 1716 1844
rect 2976 1816 3004 1856
rect 3970 1844 3976 1896
rect 4028 1884 4034 1896
rect 9122 1884 9128 1896
rect 4028 1856 9128 1884
rect 4028 1844 4034 1856
rect 9122 1844 9128 1856
rect 9180 1844 9186 1896
rect 8938 1816 8944 1828
rect 1688 1788 2774 1816
rect 2976 1788 8944 1816
rect 2746 1680 2774 1788
rect 8938 1776 8944 1788
rect 8996 1776 9002 1828
rect 6546 1680 6552 1692
rect 2746 1652 6552 1680
rect 6546 1640 6552 1652
rect 6604 1640 6610 1692
<< via1 >>
rect 3388 9766 3440 9818
rect 3452 9766 3504 9818
rect 3516 9766 3568 9818
rect 3580 9766 3632 9818
rect 3644 9766 3696 9818
rect 5826 9766 5878 9818
rect 5890 9766 5942 9818
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 8264 9766 8316 9818
rect 8328 9766 8380 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 10702 9766 10754 9818
rect 10766 9766 10818 9818
rect 10830 9766 10882 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 9956 9664 10008 9716
rect 10508 9664 10560 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 1860 9528 1912 9580
rect 1952 9460 2004 9512
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9404 9528 9456 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 9220 9392 9272 9444
rect 940 9324 992 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 1492 9163 1544 9172
rect 1492 9129 1501 9163
rect 1501 9129 1535 9163
rect 1535 9129 1544 9163
rect 1492 9120 1544 9129
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 10048 9120 10100 9172
rect 10232 9163 10284 9172
rect 10232 9129 10241 9163
rect 10241 9129 10275 9163
rect 10275 9129 10284 9163
rect 10232 9120 10284 9129
rect 10140 9052 10192 9104
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 4252 8916 4304 8968
rect 4528 8848 4580 8900
rect 2872 8780 2924 8832
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 3388 8678 3440 8730
rect 3452 8678 3504 8730
rect 3516 8678 3568 8730
rect 3580 8678 3632 8730
rect 3644 8678 3696 8730
rect 5826 8678 5878 8730
rect 5890 8678 5942 8730
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 8264 8678 8316 8730
rect 8328 8678 8380 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 10702 8678 10754 8730
rect 10766 8678 10818 8730
rect 10830 8678 10882 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 9312 8576 9364 8628
rect 10600 8508 10652 8560
rect 2044 8440 2096 8492
rect 3884 8440 3936 8492
rect 2780 8372 2832 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 9864 8440 9916 8492
rect 10508 8236 10560 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 9864 8032 9916 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 7472 7828 7524 7880
rect 8944 7828 8996 7880
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 3388 7590 3440 7642
rect 3452 7590 3504 7642
rect 3516 7590 3568 7642
rect 3580 7590 3632 7642
rect 3644 7590 3696 7642
rect 5826 7590 5878 7642
rect 5890 7590 5942 7642
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 8264 7590 8316 7642
rect 8328 7590 8380 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 10702 7590 10754 7642
rect 10766 7590 10818 7642
rect 10830 7590 10882 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 10232 7488 10284 7540
rect 9312 7420 9364 7472
rect 2596 7352 2648 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10508 7284 10560 7336
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 6828 7148 6880 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 10416 7148 10468 7157
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 9312 6876 9364 6928
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 7840 6672 7892 6724
rect 9956 6740 10008 6792
rect 10876 6740 10928 6792
rect 8760 6604 8812 6656
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 10140 6604 10192 6656
rect 3388 6502 3440 6554
rect 3452 6502 3504 6554
rect 3516 6502 3568 6554
rect 3580 6502 3632 6554
rect 3644 6502 3696 6554
rect 5826 6502 5878 6554
rect 5890 6502 5942 6554
rect 5954 6502 6006 6554
rect 6018 6502 6070 6554
rect 6082 6502 6134 6554
rect 8264 6502 8316 6554
rect 8328 6502 8380 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 10702 6502 10754 6554
rect 10766 6502 10818 6554
rect 10830 6502 10882 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 5540 6264 5592 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7840 6443 7892 6452
rect 7840 6409 7849 6443
rect 7849 6409 7883 6443
rect 7883 6409 7892 6443
rect 7840 6400 7892 6409
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 10232 6400 10284 6452
rect 8116 6264 8168 6316
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 8484 6196 8536 6248
rect 9036 6332 9088 6384
rect 8760 6264 8812 6316
rect 9864 6264 9916 6316
rect 10140 6264 10192 6316
rect 9220 6196 9272 6248
rect 940 6060 992 6112
rect 7840 6060 7892 6112
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 6828 5856 6880 5908
rect 8392 5856 8444 5908
rect 9956 5856 10008 5908
rect 6736 5720 6788 5772
rect 6184 5584 6236 5636
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 8760 5652 8812 5704
rect 7196 5584 7248 5636
rect 10048 5627 10100 5636
rect 10048 5593 10057 5627
rect 10057 5593 10091 5627
rect 10091 5593 10100 5627
rect 10048 5584 10100 5593
rect 6920 5516 6972 5568
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 8944 5516 8996 5568
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 3388 5414 3440 5466
rect 3452 5414 3504 5466
rect 3516 5414 3568 5466
rect 3580 5414 3632 5466
rect 3644 5414 3696 5466
rect 5826 5414 5878 5466
rect 5890 5414 5942 5466
rect 5954 5414 6006 5466
rect 6018 5414 6070 5466
rect 6082 5414 6134 5466
rect 8264 5414 8316 5466
rect 8328 5414 8380 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 10702 5414 10754 5466
rect 10766 5414 10818 5466
rect 10830 5414 10882 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 1768 5312 1820 5364
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 1676 5108 1728 5160
rect 4160 5176 4212 5228
rect 5448 5312 5500 5364
rect 9036 5312 9088 5364
rect 10416 5312 10468 5364
rect 6828 5244 6880 5296
rect 9312 5244 9364 5296
rect 9036 5176 9088 5228
rect 4344 5108 4396 5160
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 8944 5151 8996 5160
rect 8944 5117 8953 5151
rect 8953 5117 8987 5151
rect 8987 5117 8996 5151
rect 8944 5108 8996 5117
rect 6828 5083 6880 5092
rect 6828 5049 6837 5083
rect 6837 5049 6871 5083
rect 6871 5049 6880 5083
rect 6828 5040 6880 5049
rect 8116 5040 8168 5092
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 9312 5108 9364 5160
rect 9404 5108 9456 5160
rect 10232 5040 10284 5092
rect 940 4972 992 5024
rect 5724 4972 5776 5024
rect 7196 4972 7248 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10324 4972 10376 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 4252 4768 4304 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 6184 4768 6236 4820
rect 7012 4700 7064 4752
rect 6920 4632 6972 4684
rect 7288 4632 7340 4684
rect 8760 4632 8812 4684
rect 1952 4564 2004 4616
rect 9036 4564 9088 4616
rect 4436 4428 4488 4480
rect 8300 4496 8352 4548
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 3388 4326 3440 4378
rect 3452 4326 3504 4378
rect 3516 4326 3568 4378
rect 3580 4326 3632 4378
rect 3644 4326 3696 4378
rect 5826 4326 5878 4378
rect 5890 4326 5942 4378
rect 5954 4326 6006 4378
rect 6018 4326 6070 4378
rect 6082 4326 6134 4378
rect 8264 4326 8316 4378
rect 8328 4326 8380 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 10702 4326 10754 4378
rect 10766 4326 10818 4378
rect 10830 4326 10882 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 1768 4224 1820 4276
rect 4896 4224 4948 4276
rect 8760 4224 8812 4276
rect 9220 4224 9272 4276
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 3148 4088 3200 4140
rect 4160 4156 4212 4208
rect 5264 4156 5316 4208
rect 9128 4156 9180 4208
rect 2688 4020 2740 4072
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 7840 4088 7892 4140
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 5356 4020 5408 4072
rect 6552 4020 6604 4072
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8668 4020 8720 4072
rect 10232 4088 10284 4140
rect 9312 4020 9364 4072
rect 940 3884 992 3936
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 2964 3884 3016 3936
rect 4068 3884 4120 3936
rect 5632 3952 5684 4004
rect 4436 3884 4488 3936
rect 5356 3884 5408 3936
rect 6736 3884 6788 3936
rect 8852 3884 8904 3936
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 1768 3680 1820 3732
rect 2504 3680 2556 3732
rect 2596 3680 2648 3732
rect 3884 3680 3936 3732
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 5540 3680 5592 3732
rect 6736 3680 6788 3732
rect 7012 3680 7064 3732
rect 848 3476 900 3528
rect 4068 3612 4120 3664
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 1952 3408 2004 3460
rect 1768 3340 1820 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 2412 3340 2464 3392
rect 3976 3544 4028 3596
rect 5632 3544 5684 3596
rect 10140 3612 10192 3664
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 3240 3383 3292 3392
rect 3240 3349 3249 3383
rect 3249 3349 3283 3383
rect 3283 3349 3292 3383
rect 3240 3340 3292 3349
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 4436 3408 4488 3460
rect 5632 3451 5684 3460
rect 5632 3417 5641 3451
rect 5641 3417 5675 3451
rect 5675 3417 5684 3451
rect 5632 3408 5684 3417
rect 5724 3451 5776 3460
rect 5724 3417 5733 3451
rect 5733 3417 5767 3451
rect 5767 3417 5776 3451
rect 5724 3408 5776 3417
rect 4620 3340 4672 3392
rect 4988 3340 5040 3392
rect 5264 3340 5316 3392
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 8116 3408 8168 3460
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 7564 3340 7616 3392
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 11060 3408 11112 3460
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 3388 3238 3440 3290
rect 3452 3238 3504 3290
rect 3516 3238 3568 3290
rect 3580 3238 3632 3290
rect 3644 3238 3696 3290
rect 5826 3238 5878 3290
rect 5890 3238 5942 3290
rect 5954 3238 6006 3290
rect 6018 3238 6070 3290
rect 6082 3238 6134 3290
rect 8264 3238 8316 3290
rect 8328 3238 8380 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 10702 3238 10754 3290
rect 10766 3238 10818 3290
rect 10830 3238 10882 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 1860 3136 1912 3188
rect 2228 3136 2280 3188
rect 3056 3136 3108 3188
rect 3332 3136 3384 3188
rect 3792 3136 3844 3188
rect 3884 3136 3936 3188
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 2412 3000 2464 3052
rect 4528 3068 4580 3120
rect 4620 3068 4672 3120
rect 5356 3068 5408 3120
rect 2964 3000 3016 3052
rect 2596 2864 2648 2916
rect 4436 3000 4488 3052
rect 5448 3000 5500 3052
rect 6460 3136 6512 3188
rect 8668 3136 8720 3188
rect 8944 3136 8996 3188
rect 9312 3136 9364 3188
rect 9404 3136 9456 3188
rect 6644 3068 6696 3120
rect 6736 3068 6788 3120
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 7564 3000 7616 3052
rect 10324 3136 10376 3188
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 9036 3000 9088 3052
rect 10416 3000 10468 3052
rect 5080 2864 5132 2916
rect 10508 2932 10560 2984
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 5264 2796 5316 2848
rect 5632 2796 5684 2848
rect 6276 2796 6328 2848
rect 9128 2796 9180 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 4344 2592 4396 2644
rect 5080 2592 5132 2644
rect 6828 2592 6880 2644
rect 6920 2592 6972 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 9404 2592 9456 2644
rect 10140 2592 10192 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 7472 2524 7524 2576
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 5632 2456 5684 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 1768 2388 1820 2440
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3792 2388 3844 2440
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 7012 2456 7064 2508
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 6920 2388 6972 2440
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 8116 2388 8168 2440
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8852 2388 8904 2440
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 1492 2295 1544 2304
rect 1492 2261 1501 2295
rect 1501 2261 1535 2295
rect 1535 2261 1544 2295
rect 1492 2252 1544 2261
rect 2780 2252 2832 2304
rect 5540 2252 5592 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 10048 2320 10100 2372
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 3388 2150 3440 2202
rect 3452 2150 3504 2202
rect 3516 2150 3568 2202
rect 3580 2150 3632 2202
rect 3644 2150 3696 2202
rect 5826 2150 5878 2202
rect 5890 2150 5942 2202
rect 5954 2150 6006 2202
rect 6018 2150 6070 2202
rect 6082 2150 6134 2202
rect 8264 2150 8316 2202
rect 8328 2150 8380 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 10702 2150 10754 2202
rect 10766 2150 10818 2202
rect 10830 2150 10882 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 1492 2048 1544 2100
rect 2964 2048 3016 2100
rect 7104 2048 7156 2100
rect 3884 1980 3936 2032
rect 8208 1980 8260 2032
rect 1676 1844 1728 1896
rect 3976 1844 4028 1896
rect 9128 1844 9180 1896
rect 8944 1776 8996 1828
rect 6552 1640 6604 1692
<< metal2 >>
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 2778 11248 2834 11257
rect 2778 11183 2834 11192
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 952 9081 980 9318
rect 1504 9178 1532 9687
rect 2792 9654 2820 11183
rect 3388 9820 3696 9829
rect 3388 9818 3394 9820
rect 3450 9818 3474 9820
rect 3530 9818 3554 9820
rect 3610 9818 3634 9820
rect 3690 9818 3696 9820
rect 3450 9766 3452 9818
rect 3632 9766 3634 9818
rect 3388 9764 3394 9766
rect 3450 9764 3474 9766
rect 3530 9764 3554 9766
rect 3610 9764 3634 9766
rect 3690 9764 3696 9766
rect 3388 9755 3696 9764
rect 5826 9820 6134 9829
rect 5826 9818 5832 9820
rect 5888 9818 5912 9820
rect 5968 9818 5992 9820
rect 6048 9818 6072 9820
rect 6128 9818 6134 9820
rect 5888 9766 5890 9818
rect 6070 9766 6072 9818
rect 5826 9764 5832 9766
rect 5888 9764 5912 9766
rect 5968 9764 5992 9766
rect 6048 9764 6072 9766
rect 6128 9764 6134 9766
rect 5826 9755 6134 9764
rect 8264 9820 8572 9829
rect 8264 9818 8270 9820
rect 8326 9818 8350 9820
rect 8406 9818 8430 9820
rect 8486 9818 8510 9820
rect 8566 9818 8572 9820
rect 8326 9766 8328 9818
rect 8508 9766 8510 9818
rect 8264 9764 8270 9766
rect 8326 9764 8350 9766
rect 8406 9764 8430 9766
rect 8486 9764 8510 9766
rect 8566 9764 8572 9766
rect 8264 9755 8572 9764
rect 9968 9722 9996 11455
rect 10506 10976 10562 10985
rect 10506 10911 10562 10920
rect 10138 10432 10194 10441
rect 10060 10390 10138 10418
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 9218 9616 9274 9625
rect 1860 9580 1912 9586
rect 9218 9551 9274 9560
rect 9312 9580 9364 9586
rect 1860 9522 1912 9528
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 938 9072 994 9081
rect 938 9007 994 9016
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 940 6112 992 6118
rect 940 6054 992 6060
rect 952 5817 980 6054
rect 938 5808 994 5817
rect 938 5743 994 5752
rect 1780 5370 1808 6258
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4729 980 4966
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 3641 980 3878
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 848 3528 900 3534
rect 848 3470 900 3476
rect 860 800 888 3470
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2689 1532 2790
rect 1490 2680 1546 2689
rect 1490 2615 1546 2624
rect 1688 2553 1716 5102
rect 1780 4282 1808 5170
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1780 3738 1808 4082
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1780 2446 1808 3334
rect 1872 3194 1900 9522
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 5914 1992 9454
rect 9232 9450 9260 9551
rect 9312 9522 9364 9528
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1964 3618 1992 4558
rect 2056 3942 2084 8434
rect 2332 8378 2360 8910
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 8424 2832 8430
rect 2332 8350 2544 8378
rect 2780 8366 2832 8372
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 4049 2268 4082
rect 2226 4040 2282 4049
rect 2226 3975 2282 3984
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2516 3738 2544 8350
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2608 3738 2636 7346
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2318 3632 2374 3641
rect 1964 3590 2084 3618
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 1504 2106 1532 2246
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 1688 1902 1716 2382
rect 1676 1896 1728 1902
rect 1964 1850 1992 3402
rect 1676 1838 1728 1844
rect 1780 1822 1992 1850
rect 1780 800 1808 1822
rect 846 0 902 800
rect 1766 0 1822 800
rect 2056 762 2084 3590
rect 2318 3567 2374 3576
rect 2332 3534 2360 3567
rect 2320 3528 2372 3534
rect 2134 3496 2190 3505
rect 2320 3470 2372 3476
rect 2134 3431 2190 3440
rect 2148 3058 2176 3431
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2240 3194 2268 3334
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2424 3058 2452 3334
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2594 2952 2650 2961
rect 2594 2887 2596 2896
rect 2648 2887 2650 2896
rect 2596 2858 2648 2864
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 2700 2650 2728 4014
rect 2792 3942 2820 8366
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2884 3618 2912 8774
rect 3388 8732 3696 8741
rect 3388 8730 3394 8732
rect 3450 8730 3474 8732
rect 3530 8730 3554 8732
rect 3610 8730 3634 8732
rect 3690 8730 3696 8732
rect 3450 8678 3452 8730
rect 3632 8678 3634 8730
rect 3388 8676 3394 8678
rect 3450 8676 3474 8678
rect 3530 8676 3554 8678
rect 3610 8676 3634 8678
rect 3690 8676 3696 8678
rect 3388 8667 3696 8676
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3388 7644 3696 7653
rect 3388 7642 3394 7644
rect 3450 7642 3474 7644
rect 3530 7642 3554 7644
rect 3610 7642 3634 7644
rect 3690 7642 3696 7644
rect 3450 7590 3452 7642
rect 3632 7590 3634 7642
rect 3388 7588 3394 7590
rect 3450 7588 3474 7590
rect 3530 7588 3554 7590
rect 3610 7588 3634 7590
rect 3690 7588 3696 7590
rect 3388 7579 3696 7588
rect 3388 6556 3696 6565
rect 3388 6554 3394 6556
rect 3450 6554 3474 6556
rect 3530 6554 3554 6556
rect 3610 6554 3634 6556
rect 3690 6554 3696 6556
rect 3450 6502 3452 6554
rect 3632 6502 3634 6554
rect 3388 6500 3394 6502
rect 3450 6500 3474 6502
rect 3530 6500 3554 6502
rect 3610 6500 3634 6502
rect 3690 6500 3696 6502
rect 3388 6491 3696 6500
rect 3388 5468 3696 5477
rect 3388 5466 3394 5468
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3690 5466 3696 5468
rect 3450 5414 3452 5466
rect 3632 5414 3634 5466
rect 3388 5412 3394 5414
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3690 5412 3696 5414
rect 3388 5403 3696 5412
rect 3388 4380 3696 4389
rect 3388 4378 3394 4380
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3690 4378 3696 4380
rect 3450 4326 3452 4378
rect 3632 4326 3634 4378
rect 3388 4324 3394 4326
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3690 4324 3696 4326
rect 3388 4315 3696 4324
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2792 3590 2912 3618
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2424 1601 2452 2382
rect 2792 2310 2820 3590
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 2774 2912 3470
rect 2976 3058 3004 3878
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3068 3194 3096 3470
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2884 2746 3004 2774
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2976 2106 3004 2746
rect 3160 2666 3188 4082
rect 3896 3738 3924 8434
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 4214 4200 5170
rect 4264 4826 4292 8910
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4356 4826 4384 5102
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4298 4476 4422
rect 4264 4270 4476 4298
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3602 4016 4014
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3670 4108 3878
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3068 2638 3188 2666
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 2410 1592 2466 1601
rect 2410 1527 2466 1536
rect 2608 870 2728 898
rect 2608 762 2636 870
rect 2700 800 2728 870
rect 2056 734 2636 762
rect 2686 0 2742 800
rect 3068 762 3096 2638
rect 3252 2530 3280 3334
rect 3388 3292 3696 3301
rect 3388 3290 3394 3292
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3690 3290 3696 3292
rect 3450 3238 3452 3290
rect 3632 3238 3634 3290
rect 3388 3236 3394 3238
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3690 3236 3696 3238
rect 3388 3227 3696 3236
rect 3804 3194 3832 3470
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3194 3924 3334
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3344 2774 3372 3130
rect 4264 2774 4292 4270
rect 4540 4154 4568 8842
rect 5826 8732 6134 8741
rect 5826 8730 5832 8732
rect 5888 8730 5912 8732
rect 5968 8730 5992 8732
rect 6048 8730 6072 8732
rect 6128 8730 6134 8732
rect 5888 8678 5890 8730
rect 6070 8678 6072 8730
rect 5826 8676 5832 8678
rect 5888 8676 5912 8678
rect 5968 8676 5992 8678
rect 6048 8676 6072 8678
rect 6128 8676 6134 8678
rect 5826 8667 6134 8676
rect 8264 8732 8572 8741
rect 8264 8730 8270 8732
rect 8326 8730 8350 8732
rect 8406 8730 8430 8732
rect 8486 8730 8510 8732
rect 8566 8730 8572 8732
rect 8326 8678 8328 8730
rect 8508 8678 8510 8730
rect 8264 8676 8270 8678
rect 8326 8676 8350 8678
rect 8406 8676 8430 8678
rect 8486 8676 8510 8678
rect 8566 8676 8572 8678
rect 8264 8667 8572 8676
rect 9324 8634 9352 9522
rect 9416 9178 9444 9522
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 10060 9178 10088 10390
rect 10138 10367 10194 10376
rect 10520 9722 10548 10911
rect 10702 9820 11010 9829
rect 10702 9818 10708 9820
rect 10764 9818 10788 9820
rect 10844 9818 10868 9820
rect 10924 9818 10948 9820
rect 11004 9818 11010 9820
rect 10764 9766 10766 9818
rect 10946 9766 10948 9818
rect 10702 9764 10708 9766
rect 10764 9764 10788 9766
rect 10844 9764 10868 9766
rect 10924 9764 10948 9766
rect 11004 9764 11010 9766
rect 10702 9755 11010 9764
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10152 9110 10180 9522
rect 10230 9344 10286 9353
rect 10230 9279 10286 9288
rect 10244 9178 10272 9279
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9876 8090 9904 8434
rect 10060 8090 10088 8910
rect 10702 8732 11010 8741
rect 10702 8730 10708 8732
rect 10764 8730 10788 8732
rect 10844 8730 10868 8732
rect 10924 8730 10948 8732
rect 11004 8730 11010 8732
rect 10764 8678 10766 8730
rect 10946 8678 10948 8730
rect 10702 8676 10708 8678
rect 10764 8676 10788 8678
rect 10844 8676 10868 8678
rect 10924 8676 10948 8678
rect 11004 8676 11010 8678
rect 10702 8667 11010 8676
rect 10600 8560 10652 8566
rect 10598 8528 10600 8537
rect 10652 8528 10654 8537
rect 10598 8463 10654 8472
rect 10508 8288 10560 8294
rect 10506 8256 10508 8265
rect 10560 8256 10562 8265
rect 10506 8191 10562 8200
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 10232 7880 10284 7886
rect 10428 7857 10456 7958
rect 10232 7822 10284 7828
rect 10414 7848 10470 7857
rect 5826 7644 6134 7653
rect 5826 7642 5832 7644
rect 5888 7642 5912 7644
rect 5968 7642 5992 7644
rect 6048 7642 6072 7644
rect 6128 7642 6134 7644
rect 5888 7590 5890 7642
rect 6070 7590 6072 7642
rect 5826 7588 5832 7590
rect 5888 7588 5912 7590
rect 5968 7588 5992 7590
rect 6048 7588 6072 7590
rect 6128 7588 6134 7590
rect 5826 7579 6134 7588
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5826 6556 6134 6565
rect 5826 6554 5832 6556
rect 5888 6554 5912 6556
rect 5968 6554 5992 6556
rect 6048 6554 6072 6556
rect 6128 6554 6134 6556
rect 5888 6502 5890 6554
rect 6070 6502 6072 6554
rect 5826 6500 5832 6502
rect 5888 6500 5912 6502
rect 5968 6500 5992 6502
rect 6048 6500 6072 6502
rect 6128 6500 6134 6502
rect 5826 6491 6134 6500
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 3344 2746 4016 2774
rect 3160 2514 3280 2530
rect 3148 2508 3280 2514
rect 3200 2502 3280 2508
rect 3148 2450 3200 2456
rect 3792 2440 3844 2446
rect 3790 2408 3792 2417
rect 3884 2440 3936 2446
rect 3844 2408 3846 2417
rect 3884 2382 3936 2388
rect 3790 2343 3846 2352
rect 3388 2204 3696 2213
rect 3388 2202 3394 2204
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3690 2202 3696 2204
rect 3450 2150 3452 2202
rect 3632 2150 3634 2202
rect 3388 2148 3394 2150
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3690 2148 3696 2150
rect 3388 2139 3696 2148
rect 3896 2038 3924 2382
rect 3884 2032 3936 2038
rect 3884 1974 3936 1980
rect 3988 1902 4016 2746
rect 4080 2746 4292 2774
rect 4356 4126 4568 4154
rect 4908 4162 4936 4218
rect 5264 4208 5316 4214
rect 4908 4156 5264 4162
rect 4908 4150 5316 4156
rect 4908 4134 5304 4150
rect 3976 1896 4028 1902
rect 3976 1838 4028 1844
rect 4080 1465 4108 2746
rect 4356 2650 4384 4126
rect 5356 4072 5408 4078
rect 5354 4040 5356 4049
rect 5408 4040 5410 4049
rect 5354 3975 5410 3984
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4448 3466 4476 3878
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 4632 3126 4660 3334
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2961 4476 2994
rect 4434 2952 4490 2961
rect 4434 2887 4490 2896
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 3528 870 3648 898
rect 3528 762 3556 870
rect 3620 800 3648 870
rect 4540 800 4568 3062
rect 5000 2990 5028 3334
rect 5170 3088 5226 3097
rect 5170 3023 5226 3032
rect 4988 2984 5040 2990
rect 5040 2932 5120 2938
rect 4988 2926 5120 2932
rect 5000 2922 5120 2926
rect 5000 2916 5132 2922
rect 5000 2910 5080 2916
rect 5080 2858 5132 2864
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 5092 2650 5120 2858
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5184 2417 5212 3023
rect 5276 2854 5304 3334
rect 5368 3126 5396 3878
rect 5460 3738 5488 5306
rect 5552 5166 5580 6258
rect 6748 5778 6776 6258
rect 6840 5914 6868 7142
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 5826 5468 6134 5477
rect 5826 5466 5832 5468
rect 5888 5466 5912 5468
rect 5968 5466 5992 5468
rect 6048 5466 6072 5468
rect 6128 5466 6134 5468
rect 5888 5414 5890 5466
rect 6070 5414 6072 5466
rect 5826 5412 5832 5414
rect 5888 5412 5912 5414
rect 5968 5412 5992 5414
rect 6048 5412 6072 5414
rect 6128 5412 6134 5414
rect 5826 5403 6134 5412
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5552 3369 5580 3674
rect 5644 3602 5672 3946
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5736 3466 5764 4966
rect 6196 4826 6224 5578
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6840 5098 6868 5238
rect 6932 5166 6960 5510
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 5826 4380 6134 4389
rect 5826 4378 5832 4380
rect 5888 4378 5912 4380
rect 5968 4378 5992 4380
rect 6048 4378 6072 4380
rect 6128 4378 6134 4380
rect 5888 4326 5890 4378
rect 6070 4326 6072 4378
rect 5826 4324 5832 4326
rect 5888 4324 5912 4326
rect 5968 4324 5992 4326
rect 6048 4324 6072 4326
rect 6128 4324 6134 4326
rect 5826 4315 6134 4324
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5170 2408 5226 2417
rect 5170 2343 5226 2352
rect 5460 800 5488 2994
rect 5644 2854 5672 3402
rect 5826 3292 6134 3301
rect 5826 3290 5832 3292
rect 5888 3290 5912 3292
rect 5968 3290 5992 3292
rect 6048 3290 6072 3292
rect 6128 3290 6134 3292
rect 5888 3238 5890 3290
rect 6070 3238 6072 3290
rect 5826 3236 5832 3238
rect 5888 3236 5912 3238
rect 5968 3236 5992 3238
rect 6048 3236 6072 3238
rect 6128 3236 6134 3238
rect 5826 3227 6134 3236
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5538 2544 5594 2553
rect 5644 2514 5672 2790
rect 5538 2479 5594 2488
rect 5632 2508 5684 2514
rect 5552 2310 5580 2479
rect 5632 2450 5684 2456
rect 6196 2446 6224 4762
rect 6932 4690 6960 5102
rect 7208 5030 7236 5578
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6274 3904 6330 3913
rect 6274 3839 6330 3848
rect 6288 2854 6316 3839
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3194 6500 3334
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6184 2440 6236 2446
rect 6460 2440 6512 2446
rect 6184 2382 6236 2388
rect 6380 2400 6460 2428
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5826 2204 6134 2213
rect 5826 2202 5832 2204
rect 5888 2202 5912 2204
rect 5968 2202 5992 2204
rect 6048 2202 6072 2204
rect 6128 2202 6134 2204
rect 5888 2150 5890 2202
rect 6070 2150 6072 2202
rect 5826 2148 5832 2150
rect 5888 2148 5912 2150
rect 5968 2148 5992 2150
rect 6048 2148 6072 2150
rect 6128 2148 6134 2150
rect 5826 2139 6134 2148
rect 6380 800 6408 2400
rect 6460 2382 6512 2388
rect 6564 1698 6592 4014
rect 6736 3936 6788 3942
rect 7024 3924 7052 4694
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7102 4176 7158 4185
rect 7300 4146 7328 4626
rect 7102 4111 7158 4120
rect 7288 4140 7340 4146
rect 7116 4078 7144 4111
rect 7288 4082 7340 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6736 3878 6788 3884
rect 6932 3896 7052 3924
rect 6748 3738 6776 3878
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6734 3632 6790 3641
rect 6734 3567 6790 3576
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 3126 6684 3334
rect 6748 3126 6776 3567
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6840 2650 6868 3470
rect 6932 2650 6960 3896
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7024 2961 7052 3674
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7010 2952 7066 2961
rect 7010 2887 7066 2896
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7392 2650 7420 2994
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2582 7512 7822
rect 8264 7644 8572 7653
rect 8264 7642 8270 7644
rect 8326 7642 8350 7644
rect 8406 7642 8430 7644
rect 8486 7642 8510 7644
rect 8566 7642 8572 7644
rect 8326 7590 8328 7642
rect 8508 7590 8510 7642
rect 8264 7588 8270 7590
rect 8326 7588 8350 7590
rect 8406 7588 8430 7590
rect 8486 7588 8510 7590
rect 8566 7588 8572 7590
rect 8264 7579 8572 7588
rect 8956 6914 8984 7822
rect 10244 7546 10272 7822
rect 10414 7783 10470 7792
rect 10702 7644 11010 7653
rect 10702 7642 10708 7644
rect 10764 7642 10788 7644
rect 10844 7642 10868 7644
rect 10924 7642 10948 7644
rect 11004 7642 11010 7644
rect 10764 7590 10766 7642
rect 10946 7590 10948 7642
rect 10702 7588 10708 7590
rect 10764 7588 10788 7590
rect 10844 7588 10868 7590
rect 10924 7588 10948 7590
rect 11004 7588 11010 7590
rect 10702 7579 11010 7588
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9324 6934 9352 7414
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 8864 6886 8984 6914
rect 9312 6928 9364 6934
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 6458 7880 6666
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 8128 6322 8156 6734
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8264 6556 8572 6565
rect 8264 6554 8270 6556
rect 8326 6554 8350 6556
rect 8406 6554 8430 6556
rect 8486 6554 8510 6556
rect 8566 6554 8572 6556
rect 8326 6502 8328 6554
rect 8508 6502 8510 6554
rect 8264 6500 8270 6502
rect 8326 6500 8350 6502
rect 8406 6500 8430 6502
rect 8486 6500 8510 6502
rect 8566 6500 8572 6502
rect 8264 6491 8572 6500
rect 8772 6322 8800 6598
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 4146 7880 6054
rect 8404 5914 8432 6190
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8496 5574 8524 6190
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8264 5468 8572 5477
rect 8264 5466 8270 5468
rect 8326 5466 8350 5468
rect 8406 5466 8430 5468
rect 8486 5466 8510 5468
rect 8566 5466 8572 5468
rect 8326 5414 8328 5466
rect 8508 5414 8510 5466
rect 8264 5412 8270 5414
rect 8326 5412 8350 5414
rect 8406 5412 8430 5414
rect 8486 5412 8510 5414
rect 8566 5412 8572 5414
rect 8264 5403 8572 5412
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8128 3466 8156 5034
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4554 8340 4966
rect 8772 4690 8800 5646
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8264 4380 8572 4389
rect 8264 4378 8270 4380
rect 8326 4378 8350 4380
rect 8406 4378 8430 4380
rect 8486 4378 8510 4380
rect 8566 4378 8572 4380
rect 8326 4326 8328 4378
rect 8508 4326 8510 4378
rect 8264 4324 8270 4326
rect 8326 4324 8350 4326
rect 8406 4324 8430 4326
rect 8486 4324 8510 4326
rect 8566 4324 8572 4326
rect 8264 4315 8572 4324
rect 8772 4282 8800 4626
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8574 3496 8630 3505
rect 8116 3460 8168 3466
rect 8574 3431 8630 3440
rect 8116 3402 8168 3408
rect 8588 3398 8616 3431
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 7576 3058 7604 3334
rect 8264 3292 8572 3301
rect 8264 3290 8270 3292
rect 8326 3290 8350 3292
rect 8406 3290 8430 3292
rect 8486 3290 8510 3292
rect 8566 3290 8572 3292
rect 8326 3238 8328 3290
rect 8508 3238 8510 3290
rect 8264 3236 8270 3238
rect 8326 3236 8350 3238
rect 8406 3236 8430 3238
rect 8486 3236 8510 3238
rect 8566 3236 8572 3238
rect 8264 3227 8572 3236
rect 8680 3194 8708 4014
rect 8864 3942 8892 6886
rect 9312 6870 9364 6876
rect 9324 6458 9352 6870
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5166 8984 5510
rect 9048 5370 9076 6326
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9034 5264 9090 5273
rect 9034 5199 9036 5208
rect 9088 5199 9090 5208
rect 9036 5170 9088 5176
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 8298 2544 8354 2553
rect 7012 2508 7064 2514
rect 8298 2479 8354 2488
rect 7012 2450 7064 2456
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6552 1692 6604 1698
rect 6552 1634 6604 1640
rect 3068 734 3556 762
rect 3606 0 3662 800
rect 4526 0 4582 800
rect 5446 0 5502 800
rect 6366 0 6422 800
rect 6932 82 6960 2382
rect 7024 649 7052 2450
rect 8312 2446 8340 2479
rect 8864 2446 8892 3470
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9048 3058 9076 4558
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9232 4282 9260 6190
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9772 5772 9824 5778
rect 9876 5760 9904 6258
rect 9968 5914 9996 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9824 5732 9904 5760
rect 9772 5714 9824 5720
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5302 9352 5510
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9784 5234 9812 5714
rect 10060 5642 10088 6598
rect 10152 6322 10180 6598
rect 10244 6458 10272 7346
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10416 7200 10468 7206
rect 10414 7168 10416 7177
rect 10468 7168 10470 7177
rect 10414 7103 10470 7112
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10416 6112 10468 6118
rect 10414 6080 10416 6089
rect 10468 6080 10470 6089
rect 10414 6015 10470 6024
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9218 4176 9274 4185
rect 9324 4162 9352 5102
rect 9274 4134 9352 4162
rect 9218 4111 9274 4120
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9232 2938 9260 4111
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9324 3194 9352 4014
rect 9416 3194 9444 5102
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 10244 4593 10272 5034
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10230 4584 10286 4593
rect 10230 4519 10286 4528
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9876 3618 9904 4422
rect 10244 4146 10272 4422
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10232 3936 10284 3942
rect 10336 3924 10364 4966
rect 10284 3896 10364 3924
rect 10232 3878 10284 3884
rect 10140 3664 10192 3670
rect 9876 3590 10088 3618
rect 10140 3606 10192 3612
rect 9588 3528 9640 3534
rect 9508 3488 9588 3516
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9508 3074 9536 3488
rect 9588 3470 9640 3476
rect 9140 2910 9260 2938
rect 9416 3046 9536 3074
rect 9140 2854 9168 2910
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9416 2650 9444 3046
rect 9862 2816 9918 2825
rect 9483 2748 9791 2757
rect 9862 2751 9918 2760
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9876 2689 9904 2751
rect 9862 2680 9918 2689
rect 9404 2644 9456 2650
rect 9862 2615 9918 2624
rect 9404 2586 9456 2592
rect 10060 2530 10088 3590
rect 10152 3126 10180 3606
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10152 2650 10180 3062
rect 10244 2774 10272 3878
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 3194 10364 3470
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10428 3058 10456 5306
rect 10520 5001 10548 7278
rect 10876 6792 10928 6798
rect 10874 6760 10876 6769
rect 10928 6760 10930 6769
rect 10874 6695 10930 6704
rect 10702 6556 11010 6565
rect 10702 6554 10708 6556
rect 10764 6554 10788 6556
rect 10844 6554 10868 6556
rect 10924 6554 10948 6556
rect 11004 6554 11010 6556
rect 10764 6502 10766 6554
rect 10946 6502 10948 6554
rect 10702 6500 10708 6502
rect 10764 6500 10788 6502
rect 10844 6500 10868 6502
rect 10924 6500 10948 6502
rect 11004 6500 11010 6502
rect 10702 6491 11010 6500
rect 10702 5468 11010 5477
rect 10702 5466 10708 5468
rect 10764 5466 10788 5468
rect 10844 5466 10868 5468
rect 10924 5466 10948 5468
rect 11004 5466 11010 5468
rect 10764 5414 10766 5466
rect 10946 5414 10948 5466
rect 10702 5412 10708 5414
rect 10764 5412 10788 5414
rect 10844 5412 10868 5414
rect 10924 5412 10948 5414
rect 11004 5412 11010 5414
rect 10702 5403 11010 5412
rect 10506 4992 10562 5001
rect 10506 4927 10562 4936
rect 10702 4380 11010 4389
rect 10702 4378 10708 4380
rect 10764 4378 10788 4380
rect 10844 4378 10868 4380
rect 10924 4378 10948 4380
rect 11004 4378 11010 4380
rect 10764 4326 10766 4378
rect 10946 4326 10948 4378
rect 10702 4324 10708 4326
rect 10764 4324 10788 4326
rect 10844 4324 10868 4326
rect 10924 4324 10948 4326
rect 11004 4324 11010 4326
rect 10702 4315 11010 4324
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10702 3292 11010 3301
rect 10702 3290 10708 3292
rect 10764 3290 10788 3292
rect 10844 3290 10868 3292
rect 10924 3290 10948 3292
rect 11004 3290 11010 3292
rect 10764 3238 10766 3290
rect 10946 3238 10948 3290
rect 10702 3236 10708 3238
rect 10764 3236 10788 3238
rect 10844 3236 10868 3238
rect 10924 3236 10948 3238
rect 11004 3236 11010 3238
rect 10702 3227 11010 3236
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10244 2746 10364 2774
rect 10336 2650 10364 2746
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 9876 2514 10088 2530
rect 9864 2508 10088 2514
rect 9916 2502 10088 2508
rect 9864 2450 9916 2456
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8116 2440 8168 2446
rect 8208 2440 8260 2446
rect 8116 2382 8168 2388
rect 8206 2408 8208 2417
rect 8300 2440 8352 2446
rect 8260 2408 8262 2417
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 2106 7144 2246
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7300 870 7420 898
rect 7300 800 7328 870
rect 7010 640 7066 649
rect 7010 575 7066 584
rect 7010 96 7066 105
rect 6932 54 7010 82
rect 7010 31 7066 40
rect 7286 0 7342 800
rect 7392 762 7420 870
rect 7576 762 7604 2382
rect 8024 2304 8076 2310
rect 8022 2272 8024 2281
rect 8076 2272 8078 2281
rect 8022 2207 8078 2216
rect 8128 2009 8156 2382
rect 8300 2382 8352 2388
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8206 2343 8262 2352
rect 8264 2204 8572 2213
rect 8264 2202 8270 2204
rect 8326 2202 8350 2204
rect 8406 2202 8430 2204
rect 8486 2202 8510 2204
rect 8566 2202 8572 2204
rect 8326 2150 8328 2202
rect 8508 2150 8510 2202
rect 8264 2148 8270 2150
rect 8326 2148 8350 2150
rect 8406 2148 8430 2150
rect 8486 2148 8510 2150
rect 8566 2148 8572 2150
rect 8264 2139 8572 2148
rect 8208 2032 8260 2038
rect 8114 2000 8170 2009
rect 8208 1974 8260 1980
rect 8114 1935 8170 1944
rect 8220 800 8248 1974
rect 8956 1834 8984 2382
rect 9140 1902 9168 2382
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 8944 1828 8996 1834
rect 8944 1770 8996 1776
rect 9126 1592 9182 1601
rect 9126 1527 9182 1536
rect 9140 800 9168 1527
rect 10060 800 10088 2314
rect 10520 1737 10548 2926
rect 10702 2204 11010 2213
rect 10702 2202 10708 2204
rect 10764 2202 10788 2204
rect 10844 2202 10868 2204
rect 10924 2202 10948 2204
rect 11004 2202 11010 2204
rect 10764 2150 10766 2202
rect 10946 2150 10948 2202
rect 10702 2148 10708 2150
rect 10764 2148 10788 2150
rect 10844 2148 10868 2150
rect 10924 2148 10948 2150
rect 11004 2148 11010 2150
rect 10702 2139 11010 2148
rect 10506 1728 10562 1737
rect 10506 1663 10562 1672
rect 11072 1193 11100 3402
rect 11058 1184 11114 1193
rect 11058 1119 11114 1128
rect 7392 734 7604 762
rect 8206 0 8262 800
rect 9126 0 9182 800
rect 10046 0 10102 800
<< via2 >>
rect 9954 11464 10010 11520
rect 2778 11192 2834 11248
rect 1490 9696 1546 9752
rect 3394 9818 3450 9820
rect 3474 9818 3530 9820
rect 3554 9818 3610 9820
rect 3634 9818 3690 9820
rect 3394 9766 3440 9818
rect 3440 9766 3450 9818
rect 3474 9766 3504 9818
rect 3504 9766 3516 9818
rect 3516 9766 3530 9818
rect 3554 9766 3568 9818
rect 3568 9766 3580 9818
rect 3580 9766 3610 9818
rect 3634 9766 3644 9818
rect 3644 9766 3690 9818
rect 3394 9764 3450 9766
rect 3474 9764 3530 9766
rect 3554 9764 3610 9766
rect 3634 9764 3690 9766
rect 5832 9818 5888 9820
rect 5912 9818 5968 9820
rect 5992 9818 6048 9820
rect 6072 9818 6128 9820
rect 5832 9766 5878 9818
rect 5878 9766 5888 9818
rect 5912 9766 5942 9818
rect 5942 9766 5954 9818
rect 5954 9766 5968 9818
rect 5992 9766 6006 9818
rect 6006 9766 6018 9818
rect 6018 9766 6048 9818
rect 6072 9766 6082 9818
rect 6082 9766 6128 9818
rect 5832 9764 5888 9766
rect 5912 9764 5968 9766
rect 5992 9764 6048 9766
rect 6072 9764 6128 9766
rect 8270 9818 8326 9820
rect 8350 9818 8406 9820
rect 8430 9818 8486 9820
rect 8510 9818 8566 9820
rect 8270 9766 8316 9818
rect 8316 9766 8326 9818
rect 8350 9766 8380 9818
rect 8380 9766 8392 9818
rect 8392 9766 8406 9818
rect 8430 9766 8444 9818
rect 8444 9766 8456 9818
rect 8456 9766 8486 9818
rect 8510 9766 8520 9818
rect 8520 9766 8566 9818
rect 8270 9764 8326 9766
rect 8350 9764 8406 9766
rect 8430 9764 8486 9766
rect 8510 9764 8566 9766
rect 10506 10920 10562 10976
rect 9218 9560 9274 9616
rect 938 9016 994 9072
rect 1490 8200 1546 8256
rect 1490 6840 1546 6896
rect 938 5752 994 5808
rect 938 4664 994 4720
rect 938 3576 994 3632
rect 1490 2624 1546 2680
rect 1674 2488 1730 2544
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2226 3984 2282 4040
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2318 3576 2374 3632
rect 2134 3440 2190 3496
rect 2594 2916 2650 2952
rect 2594 2896 2596 2916
rect 2596 2896 2648 2916
rect 2648 2896 2650 2916
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 3394 8730 3450 8732
rect 3474 8730 3530 8732
rect 3554 8730 3610 8732
rect 3634 8730 3690 8732
rect 3394 8678 3440 8730
rect 3440 8678 3450 8730
rect 3474 8678 3504 8730
rect 3504 8678 3516 8730
rect 3516 8678 3530 8730
rect 3554 8678 3568 8730
rect 3568 8678 3580 8730
rect 3580 8678 3610 8730
rect 3634 8678 3644 8730
rect 3644 8678 3690 8730
rect 3394 8676 3450 8678
rect 3474 8676 3530 8678
rect 3554 8676 3610 8678
rect 3634 8676 3690 8678
rect 3394 7642 3450 7644
rect 3474 7642 3530 7644
rect 3554 7642 3610 7644
rect 3634 7642 3690 7644
rect 3394 7590 3440 7642
rect 3440 7590 3450 7642
rect 3474 7590 3504 7642
rect 3504 7590 3516 7642
rect 3516 7590 3530 7642
rect 3554 7590 3568 7642
rect 3568 7590 3580 7642
rect 3580 7590 3610 7642
rect 3634 7590 3644 7642
rect 3644 7590 3690 7642
rect 3394 7588 3450 7590
rect 3474 7588 3530 7590
rect 3554 7588 3610 7590
rect 3634 7588 3690 7590
rect 3394 6554 3450 6556
rect 3474 6554 3530 6556
rect 3554 6554 3610 6556
rect 3634 6554 3690 6556
rect 3394 6502 3440 6554
rect 3440 6502 3450 6554
rect 3474 6502 3504 6554
rect 3504 6502 3516 6554
rect 3516 6502 3530 6554
rect 3554 6502 3568 6554
rect 3568 6502 3580 6554
rect 3580 6502 3610 6554
rect 3634 6502 3644 6554
rect 3644 6502 3690 6554
rect 3394 6500 3450 6502
rect 3474 6500 3530 6502
rect 3554 6500 3610 6502
rect 3634 6500 3690 6502
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3440 5466
rect 3440 5414 3450 5466
rect 3474 5414 3504 5466
rect 3504 5414 3516 5466
rect 3516 5414 3530 5466
rect 3554 5414 3568 5466
rect 3568 5414 3580 5466
rect 3580 5414 3610 5466
rect 3634 5414 3644 5466
rect 3644 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3440 4378
rect 3440 4326 3450 4378
rect 3474 4326 3504 4378
rect 3504 4326 3516 4378
rect 3516 4326 3530 4378
rect 3554 4326 3568 4378
rect 3568 4326 3580 4378
rect 3580 4326 3610 4378
rect 3634 4326 3644 4378
rect 3644 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 2410 1536 2466 1592
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3440 3290
rect 3440 3238 3450 3290
rect 3474 3238 3504 3290
rect 3504 3238 3516 3290
rect 3516 3238 3530 3290
rect 3554 3238 3568 3290
rect 3568 3238 3580 3290
rect 3580 3238 3610 3290
rect 3634 3238 3644 3290
rect 3644 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 5832 8730 5888 8732
rect 5912 8730 5968 8732
rect 5992 8730 6048 8732
rect 6072 8730 6128 8732
rect 5832 8678 5878 8730
rect 5878 8678 5888 8730
rect 5912 8678 5942 8730
rect 5942 8678 5954 8730
rect 5954 8678 5968 8730
rect 5992 8678 6006 8730
rect 6006 8678 6018 8730
rect 6018 8678 6048 8730
rect 6072 8678 6082 8730
rect 6082 8678 6128 8730
rect 5832 8676 5888 8678
rect 5912 8676 5968 8678
rect 5992 8676 6048 8678
rect 6072 8676 6128 8678
rect 8270 8730 8326 8732
rect 8350 8730 8406 8732
rect 8430 8730 8486 8732
rect 8510 8730 8566 8732
rect 8270 8678 8316 8730
rect 8316 8678 8326 8730
rect 8350 8678 8380 8730
rect 8380 8678 8392 8730
rect 8392 8678 8406 8730
rect 8430 8678 8444 8730
rect 8444 8678 8456 8730
rect 8456 8678 8486 8730
rect 8510 8678 8520 8730
rect 8520 8678 8566 8730
rect 8270 8676 8326 8678
rect 8350 8676 8406 8678
rect 8430 8676 8486 8678
rect 8510 8676 8566 8678
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10138 10376 10194 10432
rect 10708 9818 10764 9820
rect 10788 9818 10844 9820
rect 10868 9818 10924 9820
rect 10948 9818 11004 9820
rect 10708 9766 10754 9818
rect 10754 9766 10764 9818
rect 10788 9766 10818 9818
rect 10818 9766 10830 9818
rect 10830 9766 10844 9818
rect 10868 9766 10882 9818
rect 10882 9766 10894 9818
rect 10894 9766 10924 9818
rect 10948 9766 10958 9818
rect 10958 9766 11004 9818
rect 10708 9764 10764 9766
rect 10788 9764 10844 9766
rect 10868 9764 10924 9766
rect 10948 9764 11004 9766
rect 10230 9288 10286 9344
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10708 8730 10764 8732
rect 10788 8730 10844 8732
rect 10868 8730 10924 8732
rect 10948 8730 11004 8732
rect 10708 8678 10754 8730
rect 10754 8678 10764 8730
rect 10788 8678 10818 8730
rect 10818 8678 10830 8730
rect 10830 8678 10844 8730
rect 10868 8678 10882 8730
rect 10882 8678 10894 8730
rect 10894 8678 10924 8730
rect 10948 8678 10958 8730
rect 10958 8678 11004 8730
rect 10708 8676 10764 8678
rect 10788 8676 10844 8678
rect 10868 8676 10924 8678
rect 10948 8676 11004 8678
rect 10598 8508 10600 8528
rect 10600 8508 10652 8528
rect 10652 8508 10654 8528
rect 10598 8472 10654 8508
rect 10506 8236 10508 8256
rect 10508 8236 10560 8256
rect 10560 8236 10562 8256
rect 10506 8200 10562 8236
rect 5832 7642 5888 7644
rect 5912 7642 5968 7644
rect 5992 7642 6048 7644
rect 6072 7642 6128 7644
rect 5832 7590 5878 7642
rect 5878 7590 5888 7642
rect 5912 7590 5942 7642
rect 5942 7590 5954 7642
rect 5954 7590 5968 7642
rect 5992 7590 6006 7642
rect 6006 7590 6018 7642
rect 6018 7590 6048 7642
rect 6072 7590 6082 7642
rect 6082 7590 6128 7642
rect 5832 7588 5888 7590
rect 5912 7588 5968 7590
rect 5992 7588 6048 7590
rect 6072 7588 6128 7590
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 5832 6554 5888 6556
rect 5912 6554 5968 6556
rect 5992 6554 6048 6556
rect 6072 6554 6128 6556
rect 5832 6502 5878 6554
rect 5878 6502 5888 6554
rect 5912 6502 5942 6554
rect 5942 6502 5954 6554
rect 5954 6502 5968 6554
rect 5992 6502 6006 6554
rect 6006 6502 6018 6554
rect 6018 6502 6048 6554
rect 6072 6502 6082 6554
rect 6082 6502 6128 6554
rect 5832 6500 5888 6502
rect 5912 6500 5968 6502
rect 5992 6500 6048 6502
rect 6072 6500 6128 6502
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 3790 2388 3792 2408
rect 3792 2388 3844 2408
rect 3844 2388 3846 2408
rect 3790 2352 3846 2388
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3440 2202
rect 3440 2150 3450 2202
rect 3474 2150 3504 2202
rect 3504 2150 3516 2202
rect 3516 2150 3530 2202
rect 3554 2150 3568 2202
rect 3568 2150 3580 2202
rect 3580 2150 3610 2202
rect 3634 2150 3644 2202
rect 3644 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 5354 4020 5356 4040
rect 5356 4020 5408 4040
rect 5408 4020 5410 4040
rect 5354 3984 5410 4020
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4434 2896 4490 2952
rect 4066 1400 4122 1456
rect 5170 3032 5226 3088
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 5832 5466 5888 5468
rect 5912 5466 5968 5468
rect 5992 5466 6048 5468
rect 6072 5466 6128 5468
rect 5832 5414 5878 5466
rect 5878 5414 5888 5466
rect 5912 5414 5942 5466
rect 5942 5414 5954 5466
rect 5954 5414 5968 5466
rect 5992 5414 6006 5466
rect 6006 5414 6018 5466
rect 6018 5414 6048 5466
rect 6072 5414 6082 5466
rect 6082 5414 6128 5466
rect 5832 5412 5888 5414
rect 5912 5412 5968 5414
rect 5992 5412 6048 5414
rect 6072 5412 6128 5414
rect 5832 4378 5888 4380
rect 5912 4378 5968 4380
rect 5992 4378 6048 4380
rect 6072 4378 6128 4380
rect 5832 4326 5878 4378
rect 5878 4326 5888 4378
rect 5912 4326 5942 4378
rect 5942 4326 5954 4378
rect 5954 4326 5968 4378
rect 5992 4326 6006 4378
rect 6006 4326 6018 4378
rect 6018 4326 6048 4378
rect 6072 4326 6082 4378
rect 6082 4326 6128 4378
rect 5832 4324 5888 4326
rect 5912 4324 5968 4326
rect 5992 4324 6048 4326
rect 6072 4324 6128 4326
rect 5538 3304 5594 3360
rect 5170 2352 5226 2408
rect 5832 3290 5888 3292
rect 5912 3290 5968 3292
rect 5992 3290 6048 3292
rect 6072 3290 6128 3292
rect 5832 3238 5878 3290
rect 5878 3238 5888 3290
rect 5912 3238 5942 3290
rect 5942 3238 5954 3290
rect 5954 3238 5968 3290
rect 5992 3238 6006 3290
rect 6006 3238 6018 3290
rect 6018 3238 6048 3290
rect 6072 3238 6082 3290
rect 6082 3238 6128 3290
rect 5832 3236 5888 3238
rect 5912 3236 5968 3238
rect 5992 3236 6048 3238
rect 6072 3236 6128 3238
rect 5538 2488 5594 2544
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 6274 3848 6330 3904
rect 5832 2202 5888 2204
rect 5912 2202 5968 2204
rect 5992 2202 6048 2204
rect 6072 2202 6128 2204
rect 5832 2150 5878 2202
rect 5878 2150 5888 2202
rect 5912 2150 5942 2202
rect 5942 2150 5954 2202
rect 5954 2150 5968 2202
rect 5992 2150 6006 2202
rect 6006 2150 6018 2202
rect 6018 2150 6048 2202
rect 6072 2150 6082 2202
rect 6082 2150 6128 2202
rect 5832 2148 5888 2150
rect 5912 2148 5968 2150
rect 5992 2148 6048 2150
rect 6072 2148 6128 2150
rect 7102 4120 7158 4176
rect 6734 3576 6790 3632
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7010 2896 7066 2952
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 8270 7642 8326 7644
rect 8350 7642 8406 7644
rect 8430 7642 8486 7644
rect 8510 7642 8566 7644
rect 8270 7590 8316 7642
rect 8316 7590 8326 7642
rect 8350 7590 8380 7642
rect 8380 7590 8392 7642
rect 8392 7590 8406 7642
rect 8430 7590 8444 7642
rect 8444 7590 8456 7642
rect 8456 7590 8486 7642
rect 8510 7590 8520 7642
rect 8520 7590 8566 7642
rect 8270 7588 8326 7590
rect 8350 7588 8406 7590
rect 8430 7588 8486 7590
rect 8510 7588 8566 7590
rect 10414 7792 10470 7848
rect 10708 7642 10764 7644
rect 10788 7642 10844 7644
rect 10868 7642 10924 7644
rect 10948 7642 11004 7644
rect 10708 7590 10754 7642
rect 10754 7590 10764 7642
rect 10788 7590 10818 7642
rect 10818 7590 10830 7642
rect 10830 7590 10844 7642
rect 10868 7590 10882 7642
rect 10882 7590 10894 7642
rect 10894 7590 10924 7642
rect 10948 7590 10958 7642
rect 10958 7590 11004 7642
rect 10708 7588 10764 7590
rect 10788 7588 10844 7590
rect 10868 7588 10924 7590
rect 10948 7588 11004 7590
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 8270 6554 8326 6556
rect 8350 6554 8406 6556
rect 8430 6554 8486 6556
rect 8510 6554 8566 6556
rect 8270 6502 8316 6554
rect 8316 6502 8326 6554
rect 8350 6502 8380 6554
rect 8380 6502 8392 6554
rect 8392 6502 8406 6554
rect 8430 6502 8444 6554
rect 8444 6502 8456 6554
rect 8456 6502 8486 6554
rect 8510 6502 8520 6554
rect 8520 6502 8566 6554
rect 8270 6500 8326 6502
rect 8350 6500 8406 6502
rect 8430 6500 8486 6502
rect 8510 6500 8566 6502
rect 8270 5466 8326 5468
rect 8350 5466 8406 5468
rect 8430 5466 8486 5468
rect 8510 5466 8566 5468
rect 8270 5414 8316 5466
rect 8316 5414 8326 5466
rect 8350 5414 8380 5466
rect 8380 5414 8392 5466
rect 8392 5414 8406 5466
rect 8430 5414 8444 5466
rect 8444 5414 8456 5466
rect 8456 5414 8486 5466
rect 8510 5414 8520 5466
rect 8520 5414 8566 5466
rect 8270 5412 8326 5414
rect 8350 5412 8406 5414
rect 8430 5412 8486 5414
rect 8510 5412 8566 5414
rect 8270 4378 8326 4380
rect 8350 4378 8406 4380
rect 8430 4378 8486 4380
rect 8510 4378 8566 4380
rect 8270 4326 8316 4378
rect 8316 4326 8326 4378
rect 8350 4326 8380 4378
rect 8380 4326 8392 4378
rect 8392 4326 8406 4378
rect 8430 4326 8444 4378
rect 8444 4326 8456 4378
rect 8456 4326 8486 4378
rect 8510 4326 8520 4378
rect 8520 4326 8566 4378
rect 8270 4324 8326 4326
rect 8350 4324 8406 4326
rect 8430 4324 8486 4326
rect 8510 4324 8566 4326
rect 8574 3440 8630 3496
rect 8270 3290 8326 3292
rect 8350 3290 8406 3292
rect 8430 3290 8486 3292
rect 8510 3290 8566 3292
rect 8270 3238 8316 3290
rect 8316 3238 8326 3290
rect 8350 3238 8380 3290
rect 8380 3238 8392 3290
rect 8392 3238 8406 3290
rect 8430 3238 8444 3290
rect 8444 3238 8456 3290
rect 8456 3238 8486 3290
rect 8510 3238 8520 3290
rect 8520 3238 8566 3290
rect 8270 3236 8326 3238
rect 8350 3236 8406 3238
rect 8430 3236 8486 3238
rect 8510 3236 8566 3238
rect 9034 5228 9090 5264
rect 9034 5208 9036 5228
rect 9036 5208 9088 5228
rect 9088 5208 9090 5228
rect 8298 2488 8354 2544
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 10414 7148 10416 7168
rect 10416 7148 10468 7168
rect 10468 7148 10470 7168
rect 10414 7112 10470 7148
rect 10414 6060 10416 6080
rect 10416 6060 10468 6080
rect 10468 6060 10470 6080
rect 10414 6024 10470 6060
rect 9218 4120 9274 4176
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 10230 4528 10286 4584
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9862 2760 9918 2816
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 9862 2624 9918 2680
rect 10874 6740 10876 6760
rect 10876 6740 10928 6760
rect 10928 6740 10930 6760
rect 10874 6704 10930 6740
rect 10708 6554 10764 6556
rect 10788 6554 10844 6556
rect 10868 6554 10924 6556
rect 10948 6554 11004 6556
rect 10708 6502 10754 6554
rect 10754 6502 10764 6554
rect 10788 6502 10818 6554
rect 10818 6502 10830 6554
rect 10830 6502 10844 6554
rect 10868 6502 10882 6554
rect 10882 6502 10894 6554
rect 10894 6502 10924 6554
rect 10948 6502 10958 6554
rect 10958 6502 11004 6554
rect 10708 6500 10764 6502
rect 10788 6500 10844 6502
rect 10868 6500 10924 6502
rect 10948 6500 11004 6502
rect 10708 5466 10764 5468
rect 10788 5466 10844 5468
rect 10868 5466 10924 5468
rect 10948 5466 11004 5468
rect 10708 5414 10754 5466
rect 10754 5414 10764 5466
rect 10788 5414 10818 5466
rect 10818 5414 10830 5466
rect 10830 5414 10844 5466
rect 10868 5414 10882 5466
rect 10882 5414 10894 5466
rect 10894 5414 10924 5466
rect 10948 5414 10958 5466
rect 10958 5414 11004 5466
rect 10708 5412 10764 5414
rect 10788 5412 10844 5414
rect 10868 5412 10924 5414
rect 10948 5412 11004 5414
rect 10506 4936 10562 4992
rect 10708 4378 10764 4380
rect 10788 4378 10844 4380
rect 10868 4378 10924 4380
rect 10948 4378 11004 4380
rect 10708 4326 10754 4378
rect 10754 4326 10764 4378
rect 10788 4326 10818 4378
rect 10818 4326 10830 4378
rect 10830 4326 10844 4378
rect 10868 4326 10882 4378
rect 10882 4326 10894 4378
rect 10894 4326 10924 4378
rect 10948 4326 10958 4378
rect 10958 4326 11004 4378
rect 10708 4324 10764 4326
rect 10788 4324 10844 4326
rect 10868 4324 10924 4326
rect 10948 4324 11004 4326
rect 10708 3290 10764 3292
rect 10788 3290 10844 3292
rect 10868 3290 10924 3292
rect 10948 3290 11004 3292
rect 10708 3238 10754 3290
rect 10754 3238 10764 3290
rect 10788 3238 10818 3290
rect 10818 3238 10830 3290
rect 10830 3238 10844 3290
rect 10868 3238 10882 3290
rect 10882 3238 10894 3290
rect 10894 3238 10924 3290
rect 10948 3238 10958 3290
rect 10958 3238 11004 3290
rect 10708 3236 10764 3238
rect 10788 3236 10844 3238
rect 10868 3236 10924 3238
rect 10948 3236 11004 3238
rect 8206 2388 8208 2408
rect 8208 2388 8260 2408
rect 8260 2388 8262 2408
rect 7010 584 7066 640
rect 7010 40 7066 96
rect 8022 2252 8024 2272
rect 8024 2252 8076 2272
rect 8076 2252 8078 2272
rect 8022 2216 8078 2252
rect 8206 2352 8262 2388
rect 8270 2202 8326 2204
rect 8350 2202 8406 2204
rect 8430 2202 8486 2204
rect 8510 2202 8566 2204
rect 8270 2150 8316 2202
rect 8316 2150 8326 2202
rect 8350 2150 8380 2202
rect 8380 2150 8392 2202
rect 8392 2150 8406 2202
rect 8430 2150 8444 2202
rect 8444 2150 8456 2202
rect 8456 2150 8486 2202
rect 8510 2150 8520 2202
rect 8520 2150 8566 2202
rect 8270 2148 8326 2150
rect 8350 2148 8406 2150
rect 8430 2148 8486 2150
rect 8510 2148 8566 2150
rect 8114 1944 8170 2000
rect 9126 1536 9182 1592
rect 10708 2202 10764 2204
rect 10788 2202 10844 2204
rect 10868 2202 10924 2204
rect 10948 2202 11004 2204
rect 10708 2150 10754 2202
rect 10754 2150 10764 2202
rect 10788 2150 10818 2202
rect 10818 2150 10830 2202
rect 10830 2150 10844 2202
rect 10868 2150 10882 2202
rect 10882 2150 10894 2202
rect 10894 2150 10924 2202
rect 10948 2150 10958 2202
rect 10958 2150 11004 2202
rect 10708 2148 10764 2150
rect 10788 2148 10844 2150
rect 10868 2148 10924 2150
rect 10948 2148 11004 2150
rect 10506 1672 10562 1728
rect 11058 1128 11114 1184
<< metal3 >>
rect 9949 11522 10015 11525
rect 11200 11522 12000 11552
rect 9949 11520 12000 11522
rect 9949 11464 9954 11520
rect 10010 11464 12000 11520
rect 9949 11462 12000 11464
rect 9949 11459 10015 11462
rect 11200 11432 12000 11462
rect 0 11250 800 11280
rect 2773 11250 2839 11253
rect 0 11248 2839 11250
rect 0 11192 2778 11248
rect 2834 11192 2839 11248
rect 0 11190 2839 11192
rect 0 11160 800 11190
rect 2773 11187 2839 11190
rect 10501 10978 10567 10981
rect 11200 10978 12000 11008
rect 10501 10976 12000 10978
rect 10501 10920 10506 10976
rect 10562 10920 12000 10976
rect 10501 10918 12000 10920
rect 10501 10915 10567 10918
rect 11200 10888 12000 10918
rect 10133 10434 10199 10437
rect 11200 10434 12000 10464
rect 10133 10432 12000 10434
rect 10133 10376 10138 10432
rect 10194 10376 12000 10432
rect 10133 10374 12000 10376
rect 10133 10371 10199 10374
rect 11200 10344 12000 10374
rect 0 10162 800 10192
rect 0 10102 1548 10162
rect 0 10072 800 10102
rect 1488 9757 1548 10102
rect 3384 9824 3700 9825
rect 3384 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3700 9824
rect 3384 9759 3700 9760
rect 5822 9824 6138 9825
rect 5822 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6138 9824
rect 5822 9759 6138 9760
rect 8260 9824 8576 9825
rect 8260 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8576 9824
rect 8260 9759 8576 9760
rect 10698 9824 11014 9825
rect 10698 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11014 9824
rect 11200 9800 12000 9920
rect 10698 9759 11014 9760
rect 1485 9752 1551 9757
rect 1485 9696 1490 9752
rect 1546 9696 1551 9752
rect 1485 9691 1551 9696
rect 11470 9690 11530 9800
rect 11102 9630 11530 9690
rect 9213 9618 9279 9621
rect 11102 9618 11162 9630
rect 9213 9616 11162 9618
rect 9213 9560 9218 9616
rect 9274 9560 11162 9616
rect 9213 9558 11162 9560
rect 9213 9555 9279 9558
rect 10225 9346 10291 9349
rect 11200 9346 12000 9376
rect 10225 9344 12000 9346
rect 10225 9288 10230 9344
rect 10286 9288 12000 9344
rect 10225 9286 12000 9288
rect 10225 9283 10291 9286
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 11200 9256 12000 9286
rect 9479 9215 9795 9216
rect 0 9074 800 9104
rect 933 9074 999 9077
rect 0 9072 999 9074
rect 0 9016 938 9072
rect 994 9016 999 9072
rect 0 9014 999 9016
rect 0 8984 800 9014
rect 933 9011 999 9014
rect 3384 8736 3700 8737
rect 3384 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3700 8736
rect 3384 8671 3700 8672
rect 5822 8736 6138 8737
rect 5822 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6138 8736
rect 5822 8671 6138 8672
rect 8260 8736 8576 8737
rect 8260 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8576 8736
rect 8260 8671 8576 8672
rect 10698 8736 11014 8737
rect 10698 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11014 8736
rect 11200 8712 12000 8832
rect 10698 8671 11014 8672
rect 10593 8530 10659 8533
rect 11286 8530 11346 8712
rect 10593 8528 11346 8530
rect 10593 8472 10598 8528
rect 10654 8472 11346 8528
rect 10593 8470 11346 8472
rect 10593 8467 10659 8470
rect 1485 8256 1551 8261
rect 1485 8200 1490 8256
rect 1546 8200 1551 8256
rect 1485 8195 1551 8200
rect 10501 8258 10567 8261
rect 11200 8258 12000 8288
rect 10501 8256 12000 8258
rect 10501 8200 10506 8256
rect 10562 8200 12000 8256
rect 10501 8198 12000 8200
rect 10501 8195 10567 8198
rect 0 7986 800 8016
rect 1488 7986 1548 8195
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 11200 8168 12000 8198
rect 9479 8127 9795 8128
rect 0 7926 1548 7986
rect 0 7896 800 7926
rect 10409 7850 10475 7853
rect 10409 7848 11162 7850
rect 10409 7792 10414 7848
rect 10470 7792 11162 7848
rect 10409 7790 11162 7792
rect 10409 7787 10475 7790
rect 11102 7748 11162 7790
rect 11102 7744 11346 7748
rect 11102 7688 12000 7744
rect 3384 7648 3700 7649
rect 3384 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3700 7648
rect 3384 7583 3700 7584
rect 5822 7648 6138 7649
rect 5822 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6138 7648
rect 5822 7583 6138 7584
rect 8260 7648 8576 7649
rect 8260 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8576 7648
rect 8260 7583 8576 7584
rect 10698 7648 11014 7649
rect 10698 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11014 7648
rect 11200 7624 12000 7688
rect 10698 7583 11014 7584
rect 10409 7170 10475 7173
rect 11200 7170 12000 7200
rect 10409 7168 12000 7170
rect 10409 7112 10414 7168
rect 10470 7112 12000 7168
rect 10409 7110 12000 7112
rect 10409 7107 10475 7110
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 11200 7080 12000 7110
rect 9479 7039 9795 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 10869 6762 10935 6765
rect 10869 6760 11162 6762
rect 10869 6704 10874 6760
rect 10930 6704 11162 6760
rect 10869 6702 11162 6704
rect 10869 6699 10935 6702
rect 11102 6660 11162 6702
rect 11102 6656 11346 6660
rect 11102 6600 12000 6656
rect 3384 6560 3700 6561
rect 3384 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3700 6560
rect 3384 6495 3700 6496
rect 5822 6560 6138 6561
rect 5822 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6138 6560
rect 5822 6495 6138 6496
rect 8260 6560 8576 6561
rect 8260 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8576 6560
rect 8260 6495 8576 6496
rect 10698 6560 11014 6561
rect 10698 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11014 6560
rect 11200 6536 12000 6600
rect 10698 6495 11014 6496
rect 10409 6082 10475 6085
rect 11200 6082 12000 6112
rect 10409 6080 12000 6082
rect 10409 6024 10414 6080
rect 10470 6024 12000 6080
rect 10409 6022 12000 6024
rect 10409 6019 10475 6022
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 11200 5992 12000 6022
rect 9479 5951 9795 5952
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 9630 5614 11162 5674
rect 3384 5472 3700 5473
rect 3384 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3700 5472
rect 3384 5407 3700 5408
rect 5822 5472 6138 5473
rect 5822 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6138 5472
rect 5822 5407 6138 5408
rect 8260 5472 8576 5473
rect 8260 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8576 5472
rect 8260 5407 8576 5408
rect 9029 5266 9095 5269
rect 9630 5266 9690 5614
rect 11102 5572 11162 5614
rect 11102 5568 11346 5572
rect 11102 5512 12000 5568
rect 10698 5472 11014 5473
rect 10698 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11014 5472
rect 11200 5448 12000 5512
rect 10698 5407 11014 5408
rect 9029 5264 9690 5266
rect 9029 5208 9034 5264
rect 9090 5208 9690 5264
rect 9029 5206 9690 5208
rect 9029 5203 9095 5206
rect 10501 4994 10567 4997
rect 11200 4994 12000 5024
rect 10501 4992 12000 4994
rect 10501 4936 10506 4992
rect 10562 4936 12000 4992
rect 10501 4934 12000 4936
rect 10501 4931 10567 4934
rect 2165 4928 2481 4929
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 11200 4904 12000 4934
rect 9479 4863 9795 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 10225 4586 10291 4589
rect 10225 4584 11162 4586
rect 10225 4528 10230 4584
rect 10286 4528 11162 4584
rect 10225 4526 11162 4528
rect 10225 4523 10291 4526
rect 11102 4484 11162 4526
rect 11102 4480 11346 4484
rect 11102 4424 12000 4480
rect 3384 4384 3700 4385
rect 3384 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3700 4384
rect 3384 4319 3700 4320
rect 5822 4384 6138 4385
rect 5822 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6138 4384
rect 5822 4319 6138 4320
rect 8260 4384 8576 4385
rect 8260 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8576 4384
rect 8260 4319 8576 4320
rect 10698 4384 11014 4385
rect 10698 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11014 4384
rect 11200 4360 12000 4424
rect 10698 4319 11014 4320
rect 7097 4178 7163 4181
rect 9213 4178 9279 4181
rect 7097 4176 9279 4178
rect 7097 4120 7102 4176
rect 7158 4120 9218 4176
rect 9274 4120 9279 4176
rect 7097 4118 9279 4120
rect 7097 4115 7163 4118
rect 9213 4115 9279 4118
rect 2221 4042 2287 4045
rect 5349 4042 5415 4045
rect 2221 4040 5274 4042
rect 2221 3984 2226 4040
rect 2282 3984 5274 4040
rect 2221 3982 5274 3984
rect 2221 3979 2287 3982
rect 5214 3906 5274 3982
rect 5349 4040 9920 4042
rect 5349 3984 5354 4040
rect 5410 3984 9920 4040
rect 5349 3982 9920 3984
rect 5349 3979 5415 3982
rect 6269 3906 6335 3909
rect 5214 3904 6335 3906
rect 5214 3848 6274 3904
rect 6330 3848 6335 3904
rect 5214 3846 6335 3848
rect 9860 3906 9920 3982
rect 11200 3906 12000 3936
rect 9860 3846 12000 3906
rect 6269 3843 6335 3846
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 11200 3816 12000 3846
rect 9479 3775 9795 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 2313 3634 2379 3637
rect 6729 3634 6795 3637
rect 2313 3632 6795 3634
rect 2313 3576 2318 3632
rect 2374 3576 6734 3632
rect 6790 3576 6795 3632
rect 2313 3574 6795 3576
rect 2313 3571 2379 3574
rect 6729 3571 6795 3574
rect 2129 3498 2195 3501
rect 8569 3498 8635 3501
rect 2129 3496 8635 3498
rect 2129 3440 2134 3496
rect 2190 3440 8574 3496
rect 8630 3440 8635 3496
rect 2129 3438 8635 3440
rect 2129 3435 2195 3438
rect 8569 3435 8635 3438
rect 5533 3362 5599 3365
rect 4110 3360 5599 3362
rect 4110 3304 5538 3360
rect 5594 3304 5599 3360
rect 4110 3302 5599 3304
rect 3384 3296 3700 3297
rect 3384 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3700 3296
rect 3384 3231 3700 3232
rect 2589 2954 2655 2957
rect 4110 2954 4170 3302
rect 5533 3299 5599 3302
rect 5822 3296 6138 3297
rect 5822 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6138 3296
rect 5822 3231 6138 3232
rect 8260 3296 8576 3297
rect 8260 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8576 3296
rect 8260 3231 8576 3232
rect 10698 3296 11014 3297
rect 10698 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11014 3296
rect 11200 3272 12000 3392
rect 10698 3231 11014 3232
rect 5165 3090 5231 3093
rect 11286 3090 11346 3272
rect 5165 3088 11346 3090
rect 5165 3032 5170 3088
rect 5226 3032 11346 3088
rect 5165 3030 11346 3032
rect 5165 3027 5231 3030
rect 2589 2952 4170 2954
rect 2589 2896 2594 2952
rect 2650 2896 4170 2952
rect 2589 2894 4170 2896
rect 4429 2954 4495 2957
rect 7005 2954 7071 2957
rect 4429 2952 7071 2954
rect 4429 2896 4434 2952
rect 4490 2896 7010 2952
rect 7066 2896 7071 2952
rect 4429 2894 7071 2896
rect 2589 2891 2655 2894
rect 4429 2891 4495 2894
rect 7005 2891 7071 2894
rect 9857 2818 9923 2821
rect 11200 2818 12000 2848
rect 9857 2816 12000 2818
rect 9857 2760 9862 2816
rect 9918 2760 12000 2816
rect 9857 2758 12000 2760
rect 9857 2755 9923 2758
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 11200 2728 12000 2758
rect 9479 2687 9795 2688
rect 1485 2682 1551 2685
rect 798 2680 1551 2682
rect 798 2624 1490 2680
rect 1546 2624 1551 2680
rect 798 2622 1551 2624
rect 798 2576 858 2622
rect 1485 2619 1551 2622
rect 9857 2680 9923 2685
rect 9857 2624 9862 2680
rect 9918 2624 9923 2680
rect 9857 2619 9923 2624
rect 0 2486 858 2576
rect 1669 2546 1735 2549
rect 5533 2546 5599 2549
rect 8293 2546 8359 2549
rect 1669 2544 5458 2546
rect 1669 2488 1674 2544
rect 1730 2488 5458 2544
rect 1669 2486 5458 2488
rect 0 2456 800 2486
rect 1669 2483 1735 2486
rect 3785 2410 3851 2413
rect 5165 2410 5231 2413
rect 3785 2408 5231 2410
rect 3785 2352 3790 2408
rect 3846 2352 5170 2408
rect 5226 2352 5231 2408
rect 3785 2350 5231 2352
rect 5398 2410 5458 2486
rect 5533 2544 8359 2546
rect 5533 2488 5538 2544
rect 5594 2488 8298 2544
rect 8354 2488 8359 2544
rect 5533 2486 8359 2488
rect 5533 2483 5599 2486
rect 8293 2483 8359 2486
rect 8201 2410 8267 2413
rect 9860 2410 9920 2619
rect 5398 2350 6378 2410
rect 3785 2347 3851 2350
rect 5165 2347 5231 2350
rect 6318 2274 6378 2350
rect 8201 2408 9920 2410
rect 8201 2352 8206 2408
rect 8262 2352 9920 2408
rect 8201 2350 9920 2352
rect 8201 2347 8267 2350
rect 8017 2274 8083 2277
rect 6318 2272 8083 2274
rect 6318 2216 8022 2272
rect 8078 2216 8083 2272
rect 6318 2214 8083 2216
rect 8017 2211 8083 2214
rect 3384 2208 3700 2209
rect 3384 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3700 2208
rect 3384 2143 3700 2144
rect 5822 2208 6138 2209
rect 5822 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6138 2208
rect 5822 2143 6138 2144
rect 8260 2208 8576 2209
rect 8260 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8576 2208
rect 8260 2143 8576 2144
rect 10698 2208 11014 2209
rect 10698 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11014 2208
rect 11200 2184 12000 2304
rect 10698 2143 11014 2144
rect 8109 2002 8175 2005
rect 11286 2002 11346 2184
rect 8109 2000 11346 2002
rect 8109 1944 8114 2000
rect 8170 1944 11346 2000
rect 8109 1942 11346 1944
rect 8109 1939 8175 1942
rect 10501 1730 10567 1733
rect 11200 1730 12000 1760
rect 10501 1728 12000 1730
rect 10501 1672 10506 1728
rect 10562 1672 12000 1728
rect 10501 1670 12000 1672
rect 10501 1667 10567 1670
rect 11200 1640 12000 1670
rect 2405 1594 2471 1597
rect 9121 1594 9187 1597
rect 2405 1592 9187 1594
rect 2405 1536 2410 1592
rect 2466 1536 9126 1592
rect 9182 1536 9187 1592
rect 2405 1534 9187 1536
rect 2405 1531 2471 1534
rect 9121 1531 9187 1534
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 11053 1186 11119 1189
rect 11200 1186 12000 1216
rect 11053 1184 12000 1186
rect 11053 1128 11058 1184
rect 11114 1128 12000 1184
rect 11053 1126 12000 1128
rect 11053 1123 11119 1126
rect 11200 1096 12000 1126
rect 7005 642 7071 645
rect 11200 642 12000 672
rect 7005 640 12000 642
rect 7005 584 7010 640
rect 7066 584 12000 640
rect 7005 582 12000 584
rect 7005 579 7071 582
rect 11200 552 12000 582
rect 7005 98 7071 101
rect 11200 98 12000 128
rect 7005 96 12000 98
rect 7005 40 7010 96
rect 7066 40 12000 96
rect 7005 38 12000 40
rect 7005 35 7071 38
rect 11200 8 12000 38
<< via3 >>
rect 3390 9820 3454 9824
rect 3390 9764 3394 9820
rect 3394 9764 3450 9820
rect 3450 9764 3454 9820
rect 3390 9760 3454 9764
rect 3470 9820 3534 9824
rect 3470 9764 3474 9820
rect 3474 9764 3530 9820
rect 3530 9764 3534 9820
rect 3470 9760 3534 9764
rect 3550 9820 3614 9824
rect 3550 9764 3554 9820
rect 3554 9764 3610 9820
rect 3610 9764 3614 9820
rect 3550 9760 3614 9764
rect 3630 9820 3694 9824
rect 3630 9764 3634 9820
rect 3634 9764 3690 9820
rect 3690 9764 3694 9820
rect 3630 9760 3694 9764
rect 5828 9820 5892 9824
rect 5828 9764 5832 9820
rect 5832 9764 5888 9820
rect 5888 9764 5892 9820
rect 5828 9760 5892 9764
rect 5908 9820 5972 9824
rect 5908 9764 5912 9820
rect 5912 9764 5968 9820
rect 5968 9764 5972 9820
rect 5908 9760 5972 9764
rect 5988 9820 6052 9824
rect 5988 9764 5992 9820
rect 5992 9764 6048 9820
rect 6048 9764 6052 9820
rect 5988 9760 6052 9764
rect 6068 9820 6132 9824
rect 6068 9764 6072 9820
rect 6072 9764 6128 9820
rect 6128 9764 6132 9820
rect 6068 9760 6132 9764
rect 8266 9820 8330 9824
rect 8266 9764 8270 9820
rect 8270 9764 8326 9820
rect 8326 9764 8330 9820
rect 8266 9760 8330 9764
rect 8346 9820 8410 9824
rect 8346 9764 8350 9820
rect 8350 9764 8406 9820
rect 8406 9764 8410 9820
rect 8346 9760 8410 9764
rect 8426 9820 8490 9824
rect 8426 9764 8430 9820
rect 8430 9764 8486 9820
rect 8486 9764 8490 9820
rect 8426 9760 8490 9764
rect 8506 9820 8570 9824
rect 8506 9764 8510 9820
rect 8510 9764 8566 9820
rect 8566 9764 8570 9820
rect 8506 9760 8570 9764
rect 10704 9820 10768 9824
rect 10704 9764 10708 9820
rect 10708 9764 10764 9820
rect 10764 9764 10768 9820
rect 10704 9760 10768 9764
rect 10784 9820 10848 9824
rect 10784 9764 10788 9820
rect 10788 9764 10844 9820
rect 10844 9764 10848 9820
rect 10784 9760 10848 9764
rect 10864 9820 10928 9824
rect 10864 9764 10868 9820
rect 10868 9764 10924 9820
rect 10924 9764 10928 9820
rect 10864 9760 10928 9764
rect 10944 9820 11008 9824
rect 10944 9764 10948 9820
rect 10948 9764 11004 9820
rect 11004 9764 11008 9820
rect 10944 9760 11008 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 3390 8732 3454 8736
rect 3390 8676 3394 8732
rect 3394 8676 3450 8732
rect 3450 8676 3454 8732
rect 3390 8672 3454 8676
rect 3470 8732 3534 8736
rect 3470 8676 3474 8732
rect 3474 8676 3530 8732
rect 3530 8676 3534 8732
rect 3470 8672 3534 8676
rect 3550 8732 3614 8736
rect 3550 8676 3554 8732
rect 3554 8676 3610 8732
rect 3610 8676 3614 8732
rect 3550 8672 3614 8676
rect 3630 8732 3694 8736
rect 3630 8676 3634 8732
rect 3634 8676 3690 8732
rect 3690 8676 3694 8732
rect 3630 8672 3694 8676
rect 5828 8732 5892 8736
rect 5828 8676 5832 8732
rect 5832 8676 5888 8732
rect 5888 8676 5892 8732
rect 5828 8672 5892 8676
rect 5908 8732 5972 8736
rect 5908 8676 5912 8732
rect 5912 8676 5968 8732
rect 5968 8676 5972 8732
rect 5908 8672 5972 8676
rect 5988 8732 6052 8736
rect 5988 8676 5992 8732
rect 5992 8676 6048 8732
rect 6048 8676 6052 8732
rect 5988 8672 6052 8676
rect 6068 8732 6132 8736
rect 6068 8676 6072 8732
rect 6072 8676 6128 8732
rect 6128 8676 6132 8732
rect 6068 8672 6132 8676
rect 8266 8732 8330 8736
rect 8266 8676 8270 8732
rect 8270 8676 8326 8732
rect 8326 8676 8330 8732
rect 8266 8672 8330 8676
rect 8346 8732 8410 8736
rect 8346 8676 8350 8732
rect 8350 8676 8406 8732
rect 8406 8676 8410 8732
rect 8346 8672 8410 8676
rect 8426 8732 8490 8736
rect 8426 8676 8430 8732
rect 8430 8676 8486 8732
rect 8486 8676 8490 8732
rect 8426 8672 8490 8676
rect 8506 8732 8570 8736
rect 8506 8676 8510 8732
rect 8510 8676 8566 8732
rect 8566 8676 8570 8732
rect 8506 8672 8570 8676
rect 10704 8732 10768 8736
rect 10704 8676 10708 8732
rect 10708 8676 10764 8732
rect 10764 8676 10768 8732
rect 10704 8672 10768 8676
rect 10784 8732 10848 8736
rect 10784 8676 10788 8732
rect 10788 8676 10844 8732
rect 10844 8676 10848 8732
rect 10784 8672 10848 8676
rect 10864 8732 10928 8736
rect 10864 8676 10868 8732
rect 10868 8676 10924 8732
rect 10924 8676 10928 8732
rect 10864 8672 10928 8676
rect 10944 8732 11008 8736
rect 10944 8676 10948 8732
rect 10948 8676 11004 8732
rect 11004 8676 11008 8732
rect 10944 8672 11008 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 3390 7644 3454 7648
rect 3390 7588 3394 7644
rect 3394 7588 3450 7644
rect 3450 7588 3454 7644
rect 3390 7584 3454 7588
rect 3470 7644 3534 7648
rect 3470 7588 3474 7644
rect 3474 7588 3530 7644
rect 3530 7588 3534 7644
rect 3470 7584 3534 7588
rect 3550 7644 3614 7648
rect 3550 7588 3554 7644
rect 3554 7588 3610 7644
rect 3610 7588 3614 7644
rect 3550 7584 3614 7588
rect 3630 7644 3694 7648
rect 3630 7588 3634 7644
rect 3634 7588 3690 7644
rect 3690 7588 3694 7644
rect 3630 7584 3694 7588
rect 5828 7644 5892 7648
rect 5828 7588 5832 7644
rect 5832 7588 5888 7644
rect 5888 7588 5892 7644
rect 5828 7584 5892 7588
rect 5908 7644 5972 7648
rect 5908 7588 5912 7644
rect 5912 7588 5968 7644
rect 5968 7588 5972 7644
rect 5908 7584 5972 7588
rect 5988 7644 6052 7648
rect 5988 7588 5992 7644
rect 5992 7588 6048 7644
rect 6048 7588 6052 7644
rect 5988 7584 6052 7588
rect 6068 7644 6132 7648
rect 6068 7588 6072 7644
rect 6072 7588 6128 7644
rect 6128 7588 6132 7644
rect 6068 7584 6132 7588
rect 8266 7644 8330 7648
rect 8266 7588 8270 7644
rect 8270 7588 8326 7644
rect 8326 7588 8330 7644
rect 8266 7584 8330 7588
rect 8346 7644 8410 7648
rect 8346 7588 8350 7644
rect 8350 7588 8406 7644
rect 8406 7588 8410 7644
rect 8346 7584 8410 7588
rect 8426 7644 8490 7648
rect 8426 7588 8430 7644
rect 8430 7588 8486 7644
rect 8486 7588 8490 7644
rect 8426 7584 8490 7588
rect 8506 7644 8570 7648
rect 8506 7588 8510 7644
rect 8510 7588 8566 7644
rect 8566 7588 8570 7644
rect 8506 7584 8570 7588
rect 10704 7644 10768 7648
rect 10704 7588 10708 7644
rect 10708 7588 10764 7644
rect 10764 7588 10768 7644
rect 10704 7584 10768 7588
rect 10784 7644 10848 7648
rect 10784 7588 10788 7644
rect 10788 7588 10844 7644
rect 10844 7588 10848 7644
rect 10784 7584 10848 7588
rect 10864 7644 10928 7648
rect 10864 7588 10868 7644
rect 10868 7588 10924 7644
rect 10924 7588 10928 7644
rect 10864 7584 10928 7588
rect 10944 7644 11008 7648
rect 10944 7588 10948 7644
rect 10948 7588 11004 7644
rect 11004 7588 11008 7644
rect 10944 7584 11008 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 3390 6556 3454 6560
rect 3390 6500 3394 6556
rect 3394 6500 3450 6556
rect 3450 6500 3454 6556
rect 3390 6496 3454 6500
rect 3470 6556 3534 6560
rect 3470 6500 3474 6556
rect 3474 6500 3530 6556
rect 3530 6500 3534 6556
rect 3470 6496 3534 6500
rect 3550 6556 3614 6560
rect 3550 6500 3554 6556
rect 3554 6500 3610 6556
rect 3610 6500 3614 6556
rect 3550 6496 3614 6500
rect 3630 6556 3694 6560
rect 3630 6500 3634 6556
rect 3634 6500 3690 6556
rect 3690 6500 3694 6556
rect 3630 6496 3694 6500
rect 5828 6556 5892 6560
rect 5828 6500 5832 6556
rect 5832 6500 5888 6556
rect 5888 6500 5892 6556
rect 5828 6496 5892 6500
rect 5908 6556 5972 6560
rect 5908 6500 5912 6556
rect 5912 6500 5968 6556
rect 5968 6500 5972 6556
rect 5908 6496 5972 6500
rect 5988 6556 6052 6560
rect 5988 6500 5992 6556
rect 5992 6500 6048 6556
rect 6048 6500 6052 6556
rect 5988 6496 6052 6500
rect 6068 6556 6132 6560
rect 6068 6500 6072 6556
rect 6072 6500 6128 6556
rect 6128 6500 6132 6556
rect 6068 6496 6132 6500
rect 8266 6556 8330 6560
rect 8266 6500 8270 6556
rect 8270 6500 8326 6556
rect 8326 6500 8330 6556
rect 8266 6496 8330 6500
rect 8346 6556 8410 6560
rect 8346 6500 8350 6556
rect 8350 6500 8406 6556
rect 8406 6500 8410 6556
rect 8346 6496 8410 6500
rect 8426 6556 8490 6560
rect 8426 6500 8430 6556
rect 8430 6500 8486 6556
rect 8486 6500 8490 6556
rect 8426 6496 8490 6500
rect 8506 6556 8570 6560
rect 8506 6500 8510 6556
rect 8510 6500 8566 6556
rect 8566 6500 8570 6556
rect 8506 6496 8570 6500
rect 10704 6556 10768 6560
rect 10704 6500 10708 6556
rect 10708 6500 10764 6556
rect 10764 6500 10768 6556
rect 10704 6496 10768 6500
rect 10784 6556 10848 6560
rect 10784 6500 10788 6556
rect 10788 6500 10844 6556
rect 10844 6500 10848 6556
rect 10784 6496 10848 6500
rect 10864 6556 10928 6560
rect 10864 6500 10868 6556
rect 10868 6500 10924 6556
rect 10924 6500 10928 6556
rect 10864 6496 10928 6500
rect 10944 6556 11008 6560
rect 10944 6500 10948 6556
rect 10948 6500 11004 6556
rect 11004 6500 11008 6556
rect 10944 6496 11008 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5828 5468 5892 5472
rect 5828 5412 5832 5468
rect 5832 5412 5888 5468
rect 5888 5412 5892 5468
rect 5828 5408 5892 5412
rect 5908 5468 5972 5472
rect 5908 5412 5912 5468
rect 5912 5412 5968 5468
rect 5968 5412 5972 5468
rect 5908 5408 5972 5412
rect 5988 5468 6052 5472
rect 5988 5412 5992 5468
rect 5992 5412 6048 5468
rect 6048 5412 6052 5468
rect 5988 5408 6052 5412
rect 6068 5468 6132 5472
rect 6068 5412 6072 5468
rect 6072 5412 6128 5468
rect 6128 5412 6132 5468
rect 6068 5408 6132 5412
rect 8266 5468 8330 5472
rect 8266 5412 8270 5468
rect 8270 5412 8326 5468
rect 8326 5412 8330 5468
rect 8266 5408 8330 5412
rect 8346 5468 8410 5472
rect 8346 5412 8350 5468
rect 8350 5412 8406 5468
rect 8406 5412 8410 5468
rect 8346 5408 8410 5412
rect 8426 5468 8490 5472
rect 8426 5412 8430 5468
rect 8430 5412 8486 5468
rect 8486 5412 8490 5468
rect 8426 5408 8490 5412
rect 8506 5468 8570 5472
rect 8506 5412 8510 5468
rect 8510 5412 8566 5468
rect 8566 5412 8570 5468
rect 8506 5408 8570 5412
rect 10704 5468 10768 5472
rect 10704 5412 10708 5468
rect 10708 5412 10764 5468
rect 10764 5412 10768 5468
rect 10704 5408 10768 5412
rect 10784 5468 10848 5472
rect 10784 5412 10788 5468
rect 10788 5412 10844 5468
rect 10844 5412 10848 5468
rect 10784 5408 10848 5412
rect 10864 5468 10928 5472
rect 10864 5412 10868 5468
rect 10868 5412 10924 5468
rect 10924 5412 10928 5468
rect 10864 5408 10928 5412
rect 10944 5468 11008 5472
rect 10944 5412 10948 5468
rect 10948 5412 11004 5468
rect 11004 5412 11008 5468
rect 10944 5408 11008 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5828 4380 5892 4384
rect 5828 4324 5832 4380
rect 5832 4324 5888 4380
rect 5888 4324 5892 4380
rect 5828 4320 5892 4324
rect 5908 4380 5972 4384
rect 5908 4324 5912 4380
rect 5912 4324 5968 4380
rect 5968 4324 5972 4380
rect 5908 4320 5972 4324
rect 5988 4380 6052 4384
rect 5988 4324 5992 4380
rect 5992 4324 6048 4380
rect 6048 4324 6052 4380
rect 5988 4320 6052 4324
rect 6068 4380 6132 4384
rect 6068 4324 6072 4380
rect 6072 4324 6128 4380
rect 6128 4324 6132 4380
rect 6068 4320 6132 4324
rect 8266 4380 8330 4384
rect 8266 4324 8270 4380
rect 8270 4324 8326 4380
rect 8326 4324 8330 4380
rect 8266 4320 8330 4324
rect 8346 4380 8410 4384
rect 8346 4324 8350 4380
rect 8350 4324 8406 4380
rect 8406 4324 8410 4380
rect 8346 4320 8410 4324
rect 8426 4380 8490 4384
rect 8426 4324 8430 4380
rect 8430 4324 8486 4380
rect 8486 4324 8490 4380
rect 8426 4320 8490 4324
rect 8506 4380 8570 4384
rect 8506 4324 8510 4380
rect 8510 4324 8566 4380
rect 8566 4324 8570 4380
rect 8506 4320 8570 4324
rect 10704 4380 10768 4384
rect 10704 4324 10708 4380
rect 10708 4324 10764 4380
rect 10764 4324 10768 4380
rect 10704 4320 10768 4324
rect 10784 4380 10848 4384
rect 10784 4324 10788 4380
rect 10788 4324 10844 4380
rect 10844 4324 10848 4380
rect 10784 4320 10848 4324
rect 10864 4380 10928 4384
rect 10864 4324 10868 4380
rect 10868 4324 10924 4380
rect 10924 4324 10928 4380
rect 10864 4320 10928 4324
rect 10944 4380 11008 4384
rect 10944 4324 10948 4380
rect 10948 4324 11004 4380
rect 11004 4324 11008 4380
rect 10944 4320 11008 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5828 3292 5892 3296
rect 5828 3236 5832 3292
rect 5832 3236 5888 3292
rect 5888 3236 5892 3292
rect 5828 3232 5892 3236
rect 5908 3292 5972 3296
rect 5908 3236 5912 3292
rect 5912 3236 5968 3292
rect 5968 3236 5972 3292
rect 5908 3232 5972 3236
rect 5988 3292 6052 3296
rect 5988 3236 5992 3292
rect 5992 3236 6048 3292
rect 6048 3236 6052 3292
rect 5988 3232 6052 3236
rect 6068 3292 6132 3296
rect 6068 3236 6072 3292
rect 6072 3236 6128 3292
rect 6128 3236 6132 3292
rect 6068 3232 6132 3236
rect 8266 3292 8330 3296
rect 8266 3236 8270 3292
rect 8270 3236 8326 3292
rect 8326 3236 8330 3292
rect 8266 3232 8330 3236
rect 8346 3292 8410 3296
rect 8346 3236 8350 3292
rect 8350 3236 8406 3292
rect 8406 3236 8410 3292
rect 8346 3232 8410 3236
rect 8426 3292 8490 3296
rect 8426 3236 8430 3292
rect 8430 3236 8486 3292
rect 8486 3236 8490 3292
rect 8426 3232 8490 3236
rect 8506 3292 8570 3296
rect 8506 3236 8510 3292
rect 8510 3236 8566 3292
rect 8566 3236 8570 3292
rect 8506 3232 8570 3236
rect 10704 3292 10768 3296
rect 10704 3236 10708 3292
rect 10708 3236 10764 3292
rect 10764 3236 10768 3292
rect 10704 3232 10768 3236
rect 10784 3292 10848 3296
rect 10784 3236 10788 3292
rect 10788 3236 10844 3292
rect 10844 3236 10848 3292
rect 10784 3232 10848 3236
rect 10864 3292 10928 3296
rect 10864 3236 10868 3292
rect 10868 3236 10924 3292
rect 10924 3236 10928 3292
rect 10864 3232 10928 3236
rect 10944 3292 11008 3296
rect 10944 3236 10948 3292
rect 10948 3236 11004 3292
rect 11004 3236 11008 3292
rect 10944 3232 11008 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5828 2204 5892 2208
rect 5828 2148 5832 2204
rect 5832 2148 5888 2204
rect 5888 2148 5892 2204
rect 5828 2144 5892 2148
rect 5908 2204 5972 2208
rect 5908 2148 5912 2204
rect 5912 2148 5968 2204
rect 5968 2148 5972 2204
rect 5908 2144 5972 2148
rect 5988 2204 6052 2208
rect 5988 2148 5992 2204
rect 5992 2148 6048 2204
rect 6048 2148 6052 2204
rect 5988 2144 6052 2148
rect 6068 2204 6132 2208
rect 6068 2148 6072 2204
rect 6072 2148 6128 2204
rect 6128 2148 6132 2204
rect 6068 2144 6132 2148
rect 8266 2204 8330 2208
rect 8266 2148 8270 2204
rect 8270 2148 8326 2204
rect 8326 2148 8330 2204
rect 8266 2144 8330 2148
rect 8346 2204 8410 2208
rect 8346 2148 8350 2204
rect 8350 2148 8406 2204
rect 8406 2148 8410 2204
rect 8346 2144 8410 2148
rect 8426 2204 8490 2208
rect 8426 2148 8430 2204
rect 8430 2148 8486 2204
rect 8486 2148 8490 2204
rect 8426 2144 8490 2148
rect 8506 2204 8570 2208
rect 8506 2148 8510 2204
rect 8510 2148 8566 2204
rect 8566 2148 8570 2204
rect 8506 2144 8570 2148
rect 10704 2204 10768 2208
rect 10704 2148 10708 2204
rect 10708 2148 10764 2204
rect 10764 2148 10768 2204
rect 10704 2144 10768 2148
rect 10784 2204 10848 2208
rect 10784 2148 10788 2204
rect 10788 2148 10844 2204
rect 10844 2148 10848 2204
rect 10784 2144 10848 2148
rect 10864 2204 10928 2208
rect 10864 2148 10868 2204
rect 10868 2148 10924 2204
rect 10924 2148 10928 2204
rect 10864 2144 10928 2148
rect 10944 2204 11008 2208
rect 10944 2148 10948 2204
rect 10948 2148 11004 2204
rect 11004 2148 11008 2204
rect 10944 2144 11008 2148
<< metal4 >>
rect 2163 9280 2483 9840
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 7104 2483 8128
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 4928 2483 5952
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 2752 2483 3776
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 3382 9824 3702 9840
rect 3382 9760 3390 9824
rect 3454 9760 3470 9824
rect 3534 9760 3550 9824
rect 3614 9760 3630 9824
rect 3694 9760 3702 9824
rect 3382 8736 3702 9760
rect 3382 8672 3390 8736
rect 3454 8672 3470 8736
rect 3534 8672 3550 8736
rect 3614 8672 3630 8736
rect 3694 8672 3702 8736
rect 3382 7648 3702 8672
rect 3382 7584 3390 7648
rect 3454 7584 3470 7648
rect 3534 7584 3550 7648
rect 3614 7584 3630 7648
rect 3694 7584 3702 7648
rect 3382 6560 3702 7584
rect 3382 6496 3390 6560
rect 3454 6496 3470 6560
rect 3534 6496 3550 6560
rect 3614 6496 3630 6560
rect 3694 6496 3702 6560
rect 3382 5472 3702 6496
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 4384 3702 5408
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3296 3702 4320
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2128 3702 2144
rect 4601 9280 4921 9840
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 7104 4921 8128
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 4928 4921 5952
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 2752 4921 3776
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5820 9824 6140 9840
rect 5820 9760 5828 9824
rect 5892 9760 5908 9824
rect 5972 9760 5988 9824
rect 6052 9760 6068 9824
rect 6132 9760 6140 9824
rect 5820 8736 6140 9760
rect 5820 8672 5828 8736
rect 5892 8672 5908 8736
rect 5972 8672 5988 8736
rect 6052 8672 6068 8736
rect 6132 8672 6140 8736
rect 5820 7648 6140 8672
rect 5820 7584 5828 7648
rect 5892 7584 5908 7648
rect 5972 7584 5988 7648
rect 6052 7584 6068 7648
rect 6132 7584 6140 7648
rect 5820 6560 6140 7584
rect 5820 6496 5828 6560
rect 5892 6496 5908 6560
rect 5972 6496 5988 6560
rect 6052 6496 6068 6560
rect 6132 6496 6140 6560
rect 5820 5472 6140 6496
rect 5820 5408 5828 5472
rect 5892 5408 5908 5472
rect 5972 5408 5988 5472
rect 6052 5408 6068 5472
rect 6132 5408 6140 5472
rect 5820 4384 6140 5408
rect 5820 4320 5828 4384
rect 5892 4320 5908 4384
rect 5972 4320 5988 4384
rect 6052 4320 6068 4384
rect 6132 4320 6140 4384
rect 5820 3296 6140 4320
rect 5820 3232 5828 3296
rect 5892 3232 5908 3296
rect 5972 3232 5988 3296
rect 6052 3232 6068 3296
rect 6132 3232 6140 3296
rect 5820 2208 6140 3232
rect 5820 2144 5828 2208
rect 5892 2144 5908 2208
rect 5972 2144 5988 2208
rect 6052 2144 6068 2208
rect 6132 2144 6140 2208
rect 5820 2128 6140 2144
rect 7039 9280 7359 9840
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 7104 7359 8128
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 4928 7359 5952
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 2752 7359 3776
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 8258 9824 8578 9840
rect 8258 9760 8266 9824
rect 8330 9760 8346 9824
rect 8410 9760 8426 9824
rect 8490 9760 8506 9824
rect 8570 9760 8578 9824
rect 8258 8736 8578 9760
rect 8258 8672 8266 8736
rect 8330 8672 8346 8736
rect 8410 8672 8426 8736
rect 8490 8672 8506 8736
rect 8570 8672 8578 8736
rect 8258 7648 8578 8672
rect 8258 7584 8266 7648
rect 8330 7584 8346 7648
rect 8410 7584 8426 7648
rect 8490 7584 8506 7648
rect 8570 7584 8578 7648
rect 8258 6560 8578 7584
rect 8258 6496 8266 6560
rect 8330 6496 8346 6560
rect 8410 6496 8426 6560
rect 8490 6496 8506 6560
rect 8570 6496 8578 6560
rect 8258 5472 8578 6496
rect 8258 5408 8266 5472
rect 8330 5408 8346 5472
rect 8410 5408 8426 5472
rect 8490 5408 8506 5472
rect 8570 5408 8578 5472
rect 8258 4384 8578 5408
rect 8258 4320 8266 4384
rect 8330 4320 8346 4384
rect 8410 4320 8426 4384
rect 8490 4320 8506 4384
rect 8570 4320 8578 4384
rect 8258 3296 8578 4320
rect 8258 3232 8266 3296
rect 8330 3232 8346 3296
rect 8410 3232 8426 3296
rect 8490 3232 8506 3296
rect 8570 3232 8578 3296
rect 8258 2208 8578 3232
rect 8258 2144 8266 2208
rect 8330 2144 8346 2208
rect 8410 2144 8426 2208
rect 8490 2144 8506 2208
rect 8570 2144 8578 2208
rect 8258 2128 8578 2144
rect 9477 9280 9797 9840
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 7104 9797 8128
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 4928 9797 5952
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 2752 9797 3776
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10696 9824 11016 9840
rect 10696 9760 10704 9824
rect 10768 9760 10784 9824
rect 10848 9760 10864 9824
rect 10928 9760 10944 9824
rect 11008 9760 11016 9824
rect 10696 8736 11016 9760
rect 10696 8672 10704 8736
rect 10768 8672 10784 8736
rect 10848 8672 10864 8736
rect 10928 8672 10944 8736
rect 11008 8672 11016 8736
rect 10696 7648 11016 8672
rect 10696 7584 10704 7648
rect 10768 7584 10784 7648
rect 10848 7584 10864 7648
rect 10928 7584 10944 7648
rect 11008 7584 11016 7648
rect 10696 6560 11016 7584
rect 10696 6496 10704 6560
rect 10768 6496 10784 6560
rect 10848 6496 10864 6560
rect 10928 6496 10944 6560
rect 11008 6496 11016 6560
rect 10696 5472 11016 6496
rect 10696 5408 10704 5472
rect 10768 5408 10784 5472
rect 10848 5408 10864 5472
rect 10928 5408 10944 5472
rect 11008 5408 11016 5472
rect 10696 4384 11016 5408
rect 10696 4320 10704 4384
rect 10768 4320 10784 4384
rect 10848 4320 10864 4384
rect 10928 4320 10944 4384
rect 11008 4320 11016 4384
rect 10696 3296 11016 4320
rect 10696 3232 10704 3296
rect 10768 3232 10784 3296
rect 10848 3232 10864 3296
rect 10928 3232 10944 3296
rect 11008 3232 11016 3296
rect 10696 2208 11016 3232
rect 10696 2144 10704 2208
rect 10768 2144 10784 2208
rect 10848 2144 10864 2208
rect 10928 2144 10944 2208
rect 11008 2144 11016 2208
rect 10696 2128 11016 2144
use sky130_fd_sc_hd__inv_2  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform -1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _039_
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform -1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform -1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform -1 0 8648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 8648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp 1688980957
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1688980957
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1688980957
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1688980957
transform -1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _065_
timestamp 1688980957
transform 1 0 6900 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _066_
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _067_
timestamp 1688980957
transform -1 0 5796 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _068_
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _069_
timestamp 1688980957
transform -1 0 8372 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _070_
timestamp 1688980957
transform 1 0 4048 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _071_
timestamp 1688980957
transform -1 0 5060 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform -1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform -1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _090_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _091_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _092_
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _093__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _093_
timestamp 1688980957
transform -1 0 10304 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _094__44
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _094_
timestamp 1688980957
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _095_
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _096_
timestamp 1688980957
transform -1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _097_
timestamp 1688980957
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _098_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _098__45
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _099_
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _100_
timestamp 1688980957
transform -1 0 10396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _101_
timestamp 1688980957
transform -1 0 10304 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _102_
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _103__46
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _103_
timestamp 1688980957
transform -1 0 5888 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _104_
timestamp 1688980957
transform 1 0 5520 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _105_
timestamp 1688980957
transform -1 0 5796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_61
timestamp 1688980957
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_6
timestamp 1688980957
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_20
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_24
timestamp 1688980957
transform 1 0 3312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_79
timestamp 1688980957
transform 1 0 8372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_101
timestamp 1688980957
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_83
timestamp 1688980957
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1688980957
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_12
timestamp 1688980957
transform 1 0 2208 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_24
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_36
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_87
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_10
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_64
timestamp 1688980957
transform 1 0 6992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_73
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_96
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_33
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_89
timestamp 1688980957
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_98
timestamp 1688980957
transform 1 0 10120 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_66
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_98
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_12
timestamp 1688980957
transform 1 0 2208 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_16
timestamp 1688980957
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 9844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 8372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform -1 0 9476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform -1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
flabel metal3 s 11200 5448 12000 5568 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 11200 5992 12000 6112 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 11200 552 12000 672 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 11200 1096 12000 1216 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 5 nsew signal input
flabel metal3 s 11200 1640 12000 1760 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 6 nsew signal input
flabel metal3 s 11200 2184 12000 2304 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 7 nsew signal input
flabel metal3 s 11200 2728 12000 2848 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 8 nsew signal input
flabel metal3 s 11200 3272 12000 3392 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 9 nsew signal input
flabel metal3 s 11200 3816 12000 3936 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 10 nsew signal input
flabel metal3 s 11200 4360 12000 4480 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 11 nsew signal input
flabel metal3 s 11200 4904 12000 5024 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 12 nsew signal input
flabel metal3 s 11200 7080 12000 7200 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 13 nsew signal tristate
flabel metal3 s 11200 7624 12000 7744 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 14 nsew signal tristate
flabel metal3 s 11200 8168 12000 8288 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 15 nsew signal tristate
flabel metal3 s 11200 8712 12000 8832 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 16 nsew signal tristate
flabel metal3 s 11200 9256 12000 9376 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 17 nsew signal tristate
flabel metal3 s 11200 9800 12000 9920 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 18 nsew signal tristate
flabel metal3 s 11200 10344 12000 10464 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 19 nsew signal tristate
flabel metal3 s 11200 10888 12000 11008 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 20 nsew signal tristate
flabel metal3 s 11200 11432 12000 11552 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 21 nsew signal tristate
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 22 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 23 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 24 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 25 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 26 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 27 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 28 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 29 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 30 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 31 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 32 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 33 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 34 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 35 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 36 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 37 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 38 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 39 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 prog_clk
port 40 nsew signal input
flabel metal3 s 11200 6536 12000 6656 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 41 nsew signal input
flabel metal3 s 11200 8 12000 128 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 42 nsew signal input
flabel metal4 s 2163 2128 2483 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 4601 2128 4921 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 7039 2128 7359 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 9477 2128 9797 9840 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 3382 2128 3702 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 5820 2128 6140 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 8258 2128 8578 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 10696 2128 11016 9840 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 5980 9248 5980 9248 0 vdd
rlabel via1 6060 9792 6060 9792 0 vss
rlabel metal1 3910 4046 3910 4046 0 _000_
rlabel metal2 3082 3332 3082 3332 0 _001_
rlabel metal1 3220 3026 3220 3026 0 _002_
rlabel metal1 5505 2584 5505 2584 0 _003_
rlabel metal1 7038 6290 7038 6290 0 _004_
rlabel metal2 7866 6562 7866 6562 0 _005_
rlabel metal1 9568 5882 9568 5882 0 _006_
rlabel metal1 10074 4556 10074 4556 0 _007_
rlabel metal1 9200 3162 9200 3162 0 _008_
rlabel metal1 9844 5270 9844 5270 0 _009_
rlabel metal2 9982 2516 9982 2516 0 _010_
rlabel metal2 10074 6120 10074 6120 0 _011_
rlabel metal1 9016 6970 9016 6970 0 _012_
rlabel metal1 9154 4080 9154 4080 0 _013_
rlabel metal1 8556 5882 8556 5882 0 _014_
rlabel metal1 8832 6290 8832 6290 0 _015_
rlabel metal1 6624 3094 6624 3094 0 _016_
rlabel metal2 4002 2315 4002 2315 0 _017_
rlabel metal1 9062 2618 9062 2618 0 _018_
rlabel metal1 10074 3128 10074 3128 0 _019_
rlabel metal2 3220 2516 3220 2516 0 _020_
rlabel metal1 4968 4250 4968 4250 0 _021_
rlabel metal1 5520 4998 5520 4998 0 _022_
rlabel metal2 3910 3264 3910 3264 0 _023_
rlabel metal2 874 2132 874 2132 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 10074 1554 10074 1554 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_
rlabel via2 9062 5219 9062 5219 0 ccff_head
rlabel via2 10442 6069 10442 6069 0 ccff_tail
rlabel metal1 5244 2414 5244 2414 0 chanx_right_in[0]
rlabel metal3 11186 1156 11186 1156 0 chanx_right_in[1]
rlabel metal3 10910 1700 10910 1700 0 chanx_right_in[2]
rlabel metal1 7314 2448 7314 2448 0 chanx_right_in[3]
rlabel metal3 9890 2516 9890 2516 0 chanx_right_in[4]
rlabel metal1 3358 2414 3358 2414 0 chanx_right_in[5]
rlabel metal1 2898 3026 2898 3026 0 chanx_right_in[6]
rlabel metal1 9246 5134 9246 5134 0 chanx_right_in[7]
rlabel metal1 10166 7310 10166 7310 0 chanx_right_in[8]
rlabel via2 10442 7157 10442 7157 0 chanx_right_out[0]
rlabel metal2 10442 7905 10442 7905 0 chanx_right_out[1]
rlabel metal1 10488 8262 10488 8262 0 chanx_right_out[2]
rlabel metal1 9890 8568 9890 8568 0 chanx_right_out[3]
rlabel metal2 10258 9231 10258 9231 0 chanx_right_out[4]
rlabel metal1 9200 9418 9200 9418 0 chanx_right_out[5]
rlabel metal1 9982 9146 9982 9146 0 chanx_right_out[6]
rlabel metal1 10488 9690 10488 9690 0 chanx_right_out[7]
rlabel metal1 9936 9690 9936 9690 0 chanx_right_out[8]
rlabel metal2 1794 1299 1794 1299 0 chany_bottom_in[0]
rlabel metal2 2714 823 2714 823 0 chany_bottom_in[1]
rlabel metal2 3634 823 3634 823 0 chany_bottom_in[2]
rlabel metal1 2530 3060 2530 3060 0 chany_bottom_in[3]
rlabel metal1 3450 3468 3450 3468 0 chany_bottom_in[4]
rlabel metal2 6394 1588 6394 1588 0 chany_bottom_in[5]
rlabel metal2 7314 823 7314 823 0 chany_bottom_in[6]
rlabel metal2 3910 2210 3910 2210 0 chany_bottom_in[7]
rlabel metal2 2438 1989 2438 1989 0 chany_bottom_in[8]
rlabel metal3 751 2516 751 2516 0 chany_bottom_out[0]
rlabel metal3 820 3604 820 3604 0 chany_bottom_out[1]
rlabel metal3 820 4692 820 4692 0 chany_bottom_out[2]
rlabel metal3 820 5780 820 5780 0 chany_bottom_out[3]
rlabel metal3 1096 6868 1096 6868 0 chany_bottom_out[4]
rlabel metal3 1096 7956 1096 7956 0 chany_bottom_out[5]
rlabel metal3 820 9044 820 9044 0 chany_bottom_out[6]
rlabel metal3 1096 10132 1096 10132 0 chany_bottom_out[7]
rlabel metal2 2806 10421 2806 10421 0 chany_bottom_out[8]
rlabel metal2 6210 5202 6210 5202 0 clknet_0_prog_clk
rlabel metal1 5014 2618 5014 2618 0 clknet_1_0__leaf_prog_clk
rlabel metal2 7314 4386 7314 4386 0 clknet_1_1__leaf_prog_clk
rlabel metal1 8740 5542 8740 5542 0 mem_bottom_track_1.DFF_0_.D
rlabel metal2 4462 2975 4462 2975 0 mem_bottom_track_1.DFF_0_.Q
rlabel metal1 1702 1836 1702 1836 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal2 2438 3196 2438 3196 0 mem_bottom_track_3.DFF_0_.Q
rlabel metal1 8372 4590 8372 4590 0 mem_right_track_0.DFF_0_.Q
rlabel metal1 9108 5678 9108 5678 0 mem_right_track_0.DFF_1_.Q
rlabel metal1 4968 5134 4968 5134 0 mem_right_track_2.DFF_0_.Q
rlabel metal1 10396 3162 10396 3162 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 1518 2006 1518 2006 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 9890 2618 9890 2618 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 2346 3553 2346 3553 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 5750 3060 5750 3060 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal1 2530 2482 2530 2482 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal1 5520 2822 5520 2822 0 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2070 3570 2070 3570 0 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 9982 4114 9982 4114 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 9062 2482 9062 2482 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 10350 2689 10350 2689 0 mux_right_track_0.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 9798 5474 9798 5474 0 mux_right_track_0.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 8602 6188 8602 6188 0 mux_right_track_2.INVTX1_0_.out
rlabel metal1 8004 3162 8004 3162 0 mux_right_track_2.INVTX1_1_.out
rlabel metal1 8970 6222 8970 6222 0 mux_right_track_2.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 9614 7446 9614 7446 0 mux_right_track_2.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 1886 2414 1886 2414 0 net1
rlabel metal2 5290 3094 5290 3094 0 net10
rlabel metal1 10396 3026 10396 3026 0 net11
rlabel metal1 1794 5746 1794 5746 0 net12
rlabel metal1 2484 3706 2484 3706 0 net13
rlabel metal2 4278 6868 4278 6868 0 net14
rlabel metal2 2806 6154 2806 6154 0 net15
rlabel via2 2622 2907 2622 2907 0 net16
rlabel metal1 3772 3706 3772 3706 0 net17
rlabel metal1 7084 2550 7084 2550 0 net18
rlabel metal2 7406 2822 7406 2822 0 net19
rlabel metal1 1610 2380 1610 2380 0 net2
rlabel metal2 5566 2397 5566 2397 0 net20
rlabel metal1 2714 2278 2714 2278 0 net21
rlabel metal1 10258 6630 10258 6630 0 net22
rlabel metal1 6992 2618 6992 2618 0 net23
rlabel metal1 3726 4148 3726 4148 0 net24
rlabel metal1 9982 6426 9982 6426 0 net25
rlabel metal1 10120 7514 10120 7514 0 net26
rlabel metal1 8510 8058 8510 8058 0 net27
rlabel metal1 9706 8398 9706 8398 0 net28
rlabel metal2 10074 8500 10074 8500 0 net29
rlabel metal2 6854 5168 6854 5168 0 net3
rlabel metal1 9384 8602 9384 8602 0 net30
rlabel metal1 9384 8874 9384 8874 0 net31
rlabel metal2 10166 9316 10166 9316 0 net32
rlabel metal2 9430 9350 9430 9350 0 net33
rlabel metal1 2024 3094 2024 3094 0 net34
rlabel metal1 1886 3706 1886 3706 0 net35
rlabel metal1 2070 4250 2070 4250 0 net36
rlabel metal1 1886 5338 1886 5338 0 net37
rlabel metal1 2668 3706 2668 3706 0 net38
rlabel metal1 1932 8466 1932 8466 0 net39
rlabel metal1 2162 8908 2162 8908 0 net4
rlabel metal1 1932 3162 1932 3162 0 net40
rlabel metal1 1886 8874 1886 8874 0 net41
rlabel metal1 2208 9486 2208 9486 0 net42
rlabel metal1 10258 5610 10258 5610 0 net43
rlabel metal1 9660 6766 9660 6766 0 net44
rlabel metal1 6348 2958 6348 2958 0 net45
rlabel metal1 5842 4046 5842 4046 0 net46
rlabel viali 8054 3502 8054 3502 0 net47
rlabel metal1 8367 3094 8367 3094 0 net48
rlabel metal1 4411 3434 4411 3434 0 net49
rlabel metal2 2162 3247 2162 3247 0 net5
rlabel metal1 8367 4182 8367 4182 0 net50
rlabel metal1 6588 4590 6588 4590 0 net51
rlabel metal2 7222 5304 7222 5304 0 net52
rlabel metal1 5075 3094 5075 3094 0 net53
rlabel metal2 2254 4063 2254 4063 0 net6
rlabel metal2 2990 2417 2990 2417 0 net7
rlabel metal2 1702 3825 1702 3825 0 net8
rlabel metal2 2714 3332 2714 3332 0 net9
rlabel metal3 2384 1428 2384 1428 0 prog_clk
rlabel metal1 10718 6766 10718 6766 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 6946 1241 6946 1241 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 12000 12000
<< end >>
