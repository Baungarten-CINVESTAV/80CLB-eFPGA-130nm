magic
tech sky130A
magscale 1 2
timestamp 1708041631
<< viali >>
rect 13737 17289 13771 17323
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 13829 17153 13863 17187
rect 1593 16949 1627 16983
rect 1869 16949 1903 16983
rect 1961 16949 1995 16983
rect 14381 16677 14415 16711
rect 1409 16541 1443 16575
rect 13737 16541 13771 16575
rect 14197 16541 14231 16575
rect 1593 16405 1627 16439
rect 13921 16405 13955 16439
rect 1593 15453 1627 15487
rect 2053 15453 2087 15487
rect 1777 15317 1811 15351
rect 1869 15317 1903 15351
rect 1409 14977 1443 15011
rect 14197 14977 14231 15011
rect 1593 14773 1627 14807
rect 14381 14773 14415 14807
rect 1409 13889 1443 13923
rect 1593 13753 1627 13787
rect 14381 13481 14415 13515
rect 1593 13277 1627 13311
rect 2053 13277 2087 13311
rect 13737 13277 13771 13311
rect 14197 13277 14231 13311
rect 1777 13141 1811 13175
rect 1869 13141 1903 13175
rect 13921 13141 13955 13175
rect 1593 12189 1627 12223
rect 1869 12189 1903 12223
rect 1777 12053 1811 12087
rect 2053 12053 2087 12087
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 14197 11713 14231 11747
rect 1593 11509 1627 11543
rect 1869 11509 1903 11543
rect 14381 11509 14415 11543
rect 14013 10761 14047 10795
rect 1409 10625 1443 10659
rect 14197 10625 14231 10659
rect 1593 10421 1627 10455
rect 14381 10217 14415 10251
rect 14197 10013 14231 10047
rect 1777 9945 1811 9979
rect 1501 9877 1535 9911
rect 10609 9129 10643 9163
rect 10793 8925 10827 8959
rect 1409 8857 1443 8891
rect 1777 8857 1811 8891
rect 9413 8585 9447 8619
rect 14105 8517 14139 8551
rect 1777 8449 1811 8483
rect 9597 8449 9631 8483
rect 1501 8313 1535 8347
rect 14381 8313 14415 8347
rect 8125 7497 8159 7531
rect 1777 7361 1811 7395
rect 8309 7361 8343 7395
rect 1501 7157 1535 7191
rect 6837 6953 6871 6987
rect 14381 6885 14415 6919
rect 1961 6749 1995 6783
rect 7021 6749 7055 6783
rect 11621 6749 11655 6783
rect 13277 6749 13311 6783
rect 13461 6749 13495 6783
rect 14197 6749 14231 6783
rect 1409 6681 1443 6715
rect 1777 6681 1811 6715
rect 2053 6613 2087 6647
rect 11713 6613 11747 6647
rect 13921 6613 13955 6647
rect 13093 6409 13127 6443
rect 14289 6409 14323 6443
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 11805 6273 11839 6307
rect 12081 6273 12115 6307
rect 12909 6273 12943 6307
rect 13829 6273 13863 6307
rect 14197 6273 14231 6307
rect 2145 6205 2179 6239
rect 12265 6205 12299 6239
rect 12725 6205 12759 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 13921 6205 13955 6239
rect 1869 6137 1903 6171
rect 11989 6137 12023 6171
rect 2605 6069 2639 6103
rect 2329 5865 2363 5899
rect 5549 5865 5583 5899
rect 11713 5865 11747 5899
rect 12817 5865 12851 5899
rect 13737 5865 13771 5899
rect 14197 5865 14231 5899
rect 13185 5729 13219 5763
rect 13553 5729 13587 5763
rect 1777 5661 1811 5695
rect 2053 5661 2087 5695
rect 2513 5661 2547 5695
rect 2973 5661 3007 5695
rect 5733 5661 5767 5695
rect 11529 5661 11563 5695
rect 12449 5661 12483 5695
rect 13369 5661 13403 5695
rect 13461 5661 13495 5695
rect 13921 5661 13955 5695
rect 14105 5661 14139 5695
rect 2145 5593 2179 5627
rect 1501 5525 1535 5559
rect 3065 5525 3099 5559
rect 11805 5525 11839 5559
rect 12909 5321 12943 5355
rect 13829 5321 13863 5355
rect 2421 5253 2455 5287
rect 10640 5253 10674 5287
rect 1777 5185 1811 5219
rect 3249 5185 3283 5219
rect 4169 5185 4203 5219
rect 11796 5185 11830 5219
rect 13001 5185 13035 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 14197 5185 14231 5219
rect 2145 5117 2179 5151
rect 2329 5117 2363 5151
rect 3433 5117 3467 5151
rect 7021 5117 7055 5151
rect 10885 5117 10919 5151
rect 11529 5117 11563 5151
rect 2881 5049 2915 5083
rect 3985 5049 4019 5083
rect 9505 5049 9539 5083
rect 1501 4981 1535 5015
rect 3709 4981 3743 5015
rect 6377 4981 6411 5015
rect 14381 4981 14415 5015
rect 1409 4777 1443 4811
rect 12633 4777 12667 4811
rect 13093 4709 13127 4743
rect 2789 4641 2823 4675
rect 3525 4641 3559 4675
rect 4629 4641 4663 4675
rect 5089 4641 5123 4675
rect 5457 4641 5491 4675
rect 2533 4573 2567 4607
rect 4353 4573 4387 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 11253 4573 11287 4607
rect 12909 4573 12943 4607
rect 14289 4573 14323 4607
rect 2881 4505 2915 4539
rect 3433 4505 3467 4539
rect 6561 4505 6595 4539
rect 11520 4505 11554 4539
rect 13185 4505 13219 4539
rect 13737 4505 13771 4539
rect 13829 4505 13863 4539
rect 3801 4437 3835 4471
rect 7849 4437 7883 4471
rect 14105 4437 14139 4471
rect 12173 4233 12207 4267
rect 3004 4165 3038 4199
rect 3709 4165 3743 4199
rect 4077 4165 4111 4199
rect 5181 4165 5215 4199
rect 13829 4165 13863 4199
rect 14197 4165 14231 4199
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 3801 4097 3835 4131
rect 5273 4097 5307 4131
rect 11805 4097 11839 4131
rect 12909 4097 12943 4131
rect 14105 4097 14139 4131
rect 3985 4029 4019 4063
rect 12817 4029 12851 4063
rect 13553 4029 13587 4063
rect 13921 4029 13955 4063
rect 3525 3961 3559 3995
rect 4537 3961 4571 3995
rect 1869 3893 1903 3927
rect 11897 3893 11931 3927
rect 13093 3893 13127 3927
rect 1501 3689 1535 3723
rect 12817 3689 12851 3723
rect 14381 3689 14415 3723
rect 11345 3621 11379 3655
rect 2973 3553 3007 3587
rect 13921 3553 13955 3587
rect 2053 3485 2087 3519
rect 2697 3485 2731 3519
rect 3985 3485 4019 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 13461 3485 13495 3519
rect 14197 3485 14231 3519
rect 1777 3417 1811 3451
rect 4261 3417 4295 3451
rect 4813 3417 4847 3451
rect 4905 3417 4939 3451
rect 5089 3417 5123 3451
rect 11704 3417 11738 3451
rect 12909 3417 12943 3451
rect 2145 3349 2179 3383
rect 2513 3349 2547 3383
rect 3617 3349 3651 3383
rect 4169 3349 4203 3383
rect 1869 3145 1903 3179
rect 2237 3145 2271 3179
rect 3065 3145 3099 3179
rect 4445 3145 4479 3179
rect 4721 3145 4755 3179
rect 12909 3145 12943 3179
rect 4353 3077 4387 3111
rect 7849 3077 7883 3111
rect 11796 3077 11830 3111
rect 1685 3009 1719 3043
rect 1961 3009 1995 3043
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 4629 3009 4663 3043
rect 4905 3009 4939 3043
rect 9597 3009 9631 3043
rect 11529 3009 11563 3043
rect 13001 3009 13035 3043
rect 13185 3009 13219 3043
rect 13737 2941 13771 2975
rect 13921 2941 13955 2975
rect 1593 2873 1627 2907
rect 13645 2873 13679 2907
rect 14105 2873 14139 2907
rect 2421 2805 2455 2839
rect 1593 2601 1627 2635
rect 2053 2601 2087 2635
rect 3525 2601 3559 2635
rect 5273 2601 5307 2635
rect 6377 2601 6411 2635
rect 7389 2601 7423 2635
rect 8953 2601 8987 2635
rect 9965 2601 9999 2635
rect 11529 2601 11563 2635
rect 12909 2601 12943 2635
rect 13553 2601 13587 2635
rect 13829 2601 13863 2635
rect 14197 2601 14231 2635
rect 2329 2533 2363 2567
rect 5181 2533 5215 2567
rect 12541 2533 12575 2567
rect 3065 2465 3099 2499
rect 3801 2465 3835 2499
rect 1685 2397 1719 2431
rect 2237 2397 2271 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 4057 2397 4091 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6561 2397 6595 2431
rect 7573 2397 7607 2431
rect 9137 2397 9171 2431
rect 10149 2397 10183 2431
rect 11713 2397 11747 2431
rect 12265 2397 12299 2431
rect 12725 2397 12759 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 13461 2397 13495 2431
rect 13729 2399 13763 2433
rect 14105 2397 14139 2431
rect 5549 2261 5583 2295
rect 12449 2261 12483 2295
rect 13369 2261 13403 2295
<< metal1 >>
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 13722 17280 13728 17332
rect 13780 17280 13786 17332
rect 1026 17212 1032 17264
rect 1084 17252 1090 17264
rect 1084 17224 1716 17252
rect 1084 17212 1090 17224
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1688 17193 1716 17224
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2774 17184 2780 17196
rect 2179 17156 2780 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 13814 17144 13820 17196
rect 13872 17144 13878 17196
rect 1578 16940 1584 16992
rect 1636 16940 1642 16992
rect 1854 16940 1860 16992
rect 1912 16940 1918 16992
rect 1946 16940 1952 16992
rect 2004 16940 2010 16992
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 1636 16748 13768 16776
rect 1636 16736 1642 16748
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 13740 16581 13768 16748
rect 14369 16711 14427 16717
rect 14369 16677 14381 16711
rect 14415 16677 14427 16711
rect 14369 16671 14427 16677
rect 14384 16584 14412 16671
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 992 16544 1409 16572
rect 992 16532 998 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16541 14243 16575
rect 14185 16535 14243 16541
rect 1578 16396 1584 16448
rect 1636 16396 1642 16448
rect 13909 16439 13967 16445
rect 13909 16405 13921 16439
rect 13955 16436 13967 16439
rect 14200 16436 14228 16535
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 13955 16408 14228 16436
rect 13955 16405 13967 16408
rect 13909 16399 13967 16405
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 1578 15444 1584 15496
rect 1636 15444 1642 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1688 15456 2053 15484
rect 1026 15376 1032 15428
rect 1084 15416 1090 15428
rect 1688 15416 1716 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 14182 15416 14188 15428
rect 1084 15388 1716 15416
rect 1780 15388 14188 15416
rect 1084 15376 1090 15388
rect 1780 15357 1808 15388
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 1765 15351 1823 15357
rect 1765 15317 1777 15351
rect 1811 15317 1823 15351
rect 1765 15311 1823 15317
rect 1854 15308 1860 15360
rect 1912 15308 1918 15360
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 992 14980 1409 15008
rect 992 14968 998 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 1762 14804 1768 14816
rect 1627 14776 1768 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 1762 14764 1768 14776
rect 1820 14764 1826 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 13722 13852 13728 13864
rect 1596 13824 13728 13852
rect 1596 13793 1624 13824
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13753 1639 13787
rect 1581 13747 1639 13753
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 14369 13515 14427 13521
rect 14369 13481 14381 13515
rect 14415 13512 14427 13515
rect 14415 13484 14872 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14844 13456 14872 13484
rect 14826 13404 14832 13456
rect 14884 13404 14890 13456
rect 1026 13336 1032 13388
rect 1084 13376 1090 13388
rect 1084 13348 2084 13376
rect 1084 13336 1090 13348
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 1854 13308 1860 13320
rect 1627 13280 1860 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 2056 13317 2084 13348
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 14185 13311 14243 13317
rect 14185 13277 14197 13311
rect 14231 13277 14243 13311
rect 14185 13271 14243 13277
rect 14200 13240 14228 13271
rect 1780 13212 14228 13240
rect 1780 13181 1808 13212
rect 1765 13175 1823 13181
rect 1765 13141 1777 13175
rect 1811 13141 1823 13175
rect 1765 13135 1823 13141
rect 1854 13132 1860 13184
rect 1912 13132 1918 13184
rect 13906 13132 13912 13184
rect 13964 13132 13970 13184
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 1854 12384 1860 12436
rect 1912 12384 1918 12436
rect 1872 12288 1900 12384
rect 1596 12260 1900 12288
rect 1596 12229 1624 12260
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 1762 12180 1768 12232
rect 1820 12220 1826 12232
rect 1857 12223 1915 12229
rect 1857 12220 1869 12223
rect 1820 12192 1869 12220
rect 1820 12180 1826 12192
rect 1857 12189 1869 12192
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 1765 12087 1823 12093
rect 1765 12084 1777 12087
rect 1728 12056 1777 12084
rect 1728 12044 1734 12056
rect 1765 12053 1777 12056
rect 1811 12053 1823 12087
rect 1765 12047 1823 12053
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 14182 12084 14188 12096
rect 2087 12056 14188 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1026 11636 1032 11688
rect 1084 11676 1090 11688
rect 1688 11676 1716 11707
rect 14182 11704 14188 11756
rect 14240 11704 14246 11756
rect 1084 11648 1716 11676
rect 1084 11636 1090 11648
rect 1578 11500 1584 11552
rect 1636 11500 1642 11552
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 14366 11500 14372 11552
rect 14424 11500 14430 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13872 10764 14013 10792
rect 13872 10752 13878 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 1397 10619 1455 10625
rect 6886 10628 14197 10656
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 6886 10452 6914 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 1627 10424 6914 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10248 14427 10251
rect 14415 10220 14872 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 14844 10192 14872 10220
rect 14826 10140 14832 10192
rect 14884 10140 14890 10192
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13964 10016 14197 10044
rect 13964 10004 13970 10016
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 1765 9979 1823 9985
rect 1765 9945 1777 9979
rect 1811 9976 1823 9979
rect 10594 9976 10600 9988
rect 1811 9948 10600 9976
rect 1811 9945 1823 9948
rect 1765 9939 1823 9945
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 10594 9120 10600 9172
rect 10652 9120 10658 9172
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 11054 8956 11060 8968
rect 10827 8928 11060 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 1762 8848 1768 8900
rect 1820 8848 1826 8900
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 1820 8588 9413 8616
rect 1820 8576 1826 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 1670 8508 1676 8560
rect 1728 8548 1734 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 1728 8520 14105 8548
rect 1728 8508 1734 8520
rect 14093 8517 14105 8520
rect 14139 8517 14151 8551
rect 14093 8511 14151 8517
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 5534 8480 5540 8492
rect 1811 8452 5540 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 9950 8480 9956 8492
rect 9631 8452 9956 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14458 8344 14464 8356
rect 14415 8316 14464 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 5592 7500 8125 7528
rect 5592 7488 5598 7500
rect 8113 7497 8125 7500
rect 8159 7497 8171 7531
rect 8113 7491 8171 7497
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 6822 7392 6828 7404
rect 1811 7364 6828 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 992 7160 1501 7188
rect 992 7148 998 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 6822 6944 6828 6996
rect 6880 6944 6886 6996
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6885 14427 6919
rect 14369 6879 14427 6885
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1636 6820 11652 6848
rect 1636 6808 1642 6820
rect 1946 6740 1952 6792
rect 2004 6740 2010 6792
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 11624 6789 11652 6820
rect 14384 6792 14412 6879
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13446 6740 13452 6792
rect 13504 6740 13510 6792
rect 14182 6740 14188 6792
rect 14240 6740 14246 6792
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1397 6715 1455 6721
rect 1397 6712 1409 6715
rect 992 6684 1409 6712
rect 992 6672 998 6684
rect 1397 6681 1409 6684
rect 1443 6681 1455 6715
rect 1397 6675 1455 6681
rect 1765 6715 1823 6721
rect 1765 6681 1777 6715
rect 1811 6712 1823 6715
rect 5534 6712 5540 6724
rect 1811 6684 5540 6712
rect 1811 6681 1823 6684
rect 1765 6675 1823 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 2038 6604 2044 6656
rect 2096 6604 2102 6656
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 13906 6604 13912 6656
rect 13964 6604 13970 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 11698 6400 11704 6452
rect 11756 6400 11762 6452
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13446 6440 13452 6452
rect 13127 6412 13452 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 14240 6412 14289 6440
rect 14240 6400 14246 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2056 6304 2084 6400
rect 11716 6372 11744 6400
rect 11716 6344 12112 6372
rect 1995 6276 2084 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 12084 6313 12112 6344
rect 13262 6332 13268 6384
rect 13320 6332 13326 6384
rect 13906 6332 13912 6384
rect 13964 6332 13970 6384
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6304 12955 6307
rect 13078 6304 13084 6316
rect 12943 6276 13084 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13280 6304 13308 6332
rect 13817 6307 13875 6313
rect 13280 6276 13492 6304
rect 2133 6239 2191 6245
rect 2133 6236 2145 6239
rect 1872 6208 2145 6236
rect 1872 6177 1900 6208
rect 2133 6205 2145 6208
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 12802 6236 12808 6248
rect 12759 6208 12808 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6137 1915 6171
rect 1857 6131 1915 6137
rect 11977 6171 12035 6177
rect 11977 6137 11989 6171
rect 12023 6168 12035 6171
rect 12268 6168 12296 6199
rect 12802 6196 12808 6208
rect 12860 6236 12866 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 12860 6208 13185 6236
rect 12860 6196 12866 6208
rect 13173 6205 13185 6208
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6205 13415 6239
rect 13464 6236 13492 6276
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 13924 6304 13952 6332
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13863 6276 14197 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13464 6208 13921 6236
rect 13357 6199 13415 6205
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 12023 6140 12296 6168
rect 13372 6168 13400 6199
rect 14182 6168 14188 6180
rect 13372 6140 14188 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 2593 6103 2651 6109
rect 2593 6069 2605 6103
rect 2639 6100 2651 6103
rect 3418 6100 3424 6112
rect 2639 6072 3424 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 1728 5868 2329 5896
rect 1728 5856 1734 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 2317 5859 2375 5865
rect 5534 5856 5540 5908
rect 5592 5856 5598 5908
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 11790 5896 11796 5908
rect 11747 5868 11796 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13320 5868 13737 5896
rect 13320 5856 13326 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 4706 5828 4712 5840
rect 1780 5800 4712 5828
rect 1780 5701 1808 5800
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 12618 5828 12624 5840
rect 11532 5800 12624 5828
rect 5534 5760 5540 5772
rect 2516 5732 5540 5760
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 2516 5701 2544 5732
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3007 5664 3832 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 3142 5624 3148 5636
rect 2179 5596 3148 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 3804 5568 3832 5664
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 11532 5701 11560 5800
rect 12618 5788 12624 5800
rect 12676 5828 12682 5840
rect 12676 5800 13676 5828
rect 12676 5788 12682 5800
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13219 5732 13553 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 13648 5704 13676 5800
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 13630 5692 13636 5704
rect 13495 5664 13636 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 3786 5516 3792 5568
rect 3844 5516 3850 5568
rect 11790 5516 11796 5568
rect 11848 5516 11854 5568
rect 12452 5556 12480 5652
rect 13372 5624 13400 5655
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5692 13967 5695
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13955 5664 14105 5692
rect 13955 5661 13967 5664
rect 13909 5655 13967 5661
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 13814 5624 13820 5636
rect 13372 5596 13820 5624
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 13924 5556 13952 5655
rect 12452 5528 13952 5556
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 11790 5312 11796 5364
rect 11848 5312 11854 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12492 5324 12909 5352
rect 12492 5312 12498 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 13814 5312 13820 5364
rect 13872 5312 13878 5364
rect 2406 5244 2412 5296
rect 2464 5244 2470 5296
rect 10628 5287 10686 5293
rect 10628 5253 10640 5287
rect 10674 5284 10686 5287
rect 11808 5284 11836 5312
rect 10674 5256 11836 5284
rect 10674 5253 10686 5256
rect 10628 5247 10686 5253
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2038 5216 2044 5228
rect 1811 5188 2044 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 3200 5188 3249 5216
rect 3200 5176 3206 5188
rect 3237 5185 3249 5188
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4246 5216 4252 5228
rect 4203 5188 4252 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 11784 5219 11842 5225
rect 11784 5185 11796 5219
rect 11830 5216 11842 5219
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 11830 5188 13001 5216
rect 11830 5185 11842 5188
rect 11784 5179 11842 5185
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5148 2191 5151
rect 2317 5151 2375 5157
rect 2317 5148 2329 5151
rect 2179 5120 2329 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 2317 5117 2329 5120
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5049 2927 5083
rect 3436 5080 3464 5111
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 5592 5120 7021 5148
rect 5592 5108 5598 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 10873 5151 10931 5157
rect 7055 5120 9536 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 9508 5089 9536 5120
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 11146 5148 11152 5160
rect 10919 5120 11152 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11146 5108 11152 5120
rect 11204 5148 11210 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11204 5120 11529 5148
rect 11204 5108 11210 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13740 5148 13768 5179
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 12768 5120 13768 5148
rect 12768 5108 12774 5120
rect 3973 5083 4031 5089
rect 3973 5080 3985 5083
rect 3436 5052 3985 5080
rect 2869 5043 2927 5049
rect 3973 5049 3985 5052
rect 4019 5049 4031 5083
rect 3973 5043 4031 5049
rect 9493 5083 9551 5089
rect 9493 5049 9505 5083
rect 9539 5049 9551 5083
rect 9493 5043 9551 5049
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2884 5012 2912 5043
rect 2372 4984 2912 5012
rect 2372 4972 2378 4984
rect 3694 4972 3700 5024
rect 3752 4972 3758 5024
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 4488 4984 6377 5012
rect 4488 4972 4494 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6365 4975 6423 4981
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 2498 4808 2504 4820
rect 1443 4780 2504 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 2498 4768 2504 4780
rect 2556 4808 2562 4820
rect 3786 4808 3792 4820
rect 2556 4780 3792 4808
rect 2556 4768 2562 4780
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4430 4768 4436 4820
rect 4488 4768 4494 4820
rect 12618 4768 12624 4820
rect 12676 4768 12682 4820
rect 4448 4740 4476 4768
rect 2884 4712 4476 4740
rect 13081 4743 13139 4749
rect 2774 4632 2780 4684
rect 2832 4632 2838 4684
rect 2521 4607 2579 4613
rect 2521 4573 2533 4607
rect 2567 4604 2579 4607
rect 2884 4604 2912 4712
rect 13081 4709 13093 4743
rect 13127 4709 13139 4743
rect 13081 4703 13139 4709
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 3513 4675 3571 4681
rect 3513 4672 3525 4675
rect 3476 4644 3525 4672
rect 3476 4632 3482 4644
rect 3513 4641 3525 4644
rect 3559 4672 3571 4675
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 3559 4644 4629 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5123 4644 5457 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 13096 4672 13124 4703
rect 13096 4644 14320 4672
rect 5445 4635 5503 4641
rect 2567 4576 2912 4604
rect 2567 4573 2579 4576
rect 2521 4567 2579 4573
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 3844 4576 4353 4604
rect 3844 4564 3850 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 5224 4576 5273 4604
rect 5224 4564 5230 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 14292 4613 14320 4644
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 9088 4576 11253 4604
rect 9088 4564 9094 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 11241 4567 11299 4573
rect 12820 4576 12909 4604
rect 1854 4496 1860 4548
rect 1912 4536 1918 4548
rect 2314 4536 2320 4548
rect 1912 4508 2320 4536
rect 1912 4496 1918 4508
rect 2314 4496 2320 4508
rect 2372 4536 2378 4548
rect 2869 4539 2927 4545
rect 2869 4536 2881 4539
rect 2372 4508 2881 4536
rect 2372 4496 2378 4508
rect 2869 4505 2881 4508
rect 2915 4505 2927 4539
rect 2869 4499 2927 4505
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 3421 4539 3479 4545
rect 3421 4536 3433 4539
rect 3108 4508 3433 4536
rect 3108 4496 3114 4508
rect 3421 4505 3433 4508
rect 3467 4505 3479 4539
rect 3421 4499 3479 4505
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 6549 4539 6607 4545
rect 6549 4536 6561 4539
rect 4212 4508 6561 4536
rect 4212 4496 4218 4508
rect 6549 4505 6561 4508
rect 6595 4505 6607 4539
rect 6549 4499 6607 4505
rect 11508 4539 11566 4545
rect 11508 4505 11520 4539
rect 11554 4536 11566 4539
rect 12158 4536 12164 4548
rect 11554 4508 12164 4536
rect 11554 4505 11566 4508
rect 11508 4499 11566 4505
rect 12158 4496 12164 4508
rect 12216 4496 12222 4548
rect 12820 4480 12848 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 13173 4539 13231 4545
rect 13173 4505 13185 4539
rect 13219 4536 13231 4539
rect 13538 4536 13544 4548
rect 13219 4508 13544 4536
rect 13219 4505 13231 4508
rect 13173 4499 13231 4505
rect 13538 4496 13544 4508
rect 13596 4496 13602 4548
rect 13725 4539 13783 4545
rect 13725 4505 13737 4539
rect 13771 4505 13783 4539
rect 13725 4499 13783 4505
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3200 4440 3801 4468
rect 3200 4428 3206 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 7837 4471 7895 4477
rect 7837 4468 7849 4471
rect 7708 4440 7849 4468
rect 7708 4428 7714 4440
rect 7837 4437 7849 4440
rect 7883 4437 7895 4471
rect 7837 4431 7895 4437
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 13740 4468 13768 4499
rect 13814 4496 13820 4548
rect 13872 4496 13878 4548
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13740 4440 14105 4468
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 9030 4264 9036 4276
rect 2832 4236 9036 4264
rect 2832 4224 2838 4236
rect 2992 4199 3050 4205
rect 2992 4165 3004 4199
rect 3038 4196 3050 4199
rect 3142 4196 3148 4208
rect 3038 4168 3148 4196
rect 3038 4165 3050 4168
rect 2992 4159 3050 4165
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 3252 4140 3280 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 12158 4224 12164 4276
rect 12216 4224 12222 4276
rect 3697 4199 3755 4205
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 4065 4199 4123 4205
rect 4065 4196 4077 4199
rect 3743 4168 4077 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 4065 4165 4077 4168
rect 4111 4165 4123 4199
rect 4065 4159 4123 4165
rect 5166 4156 5172 4208
rect 5224 4156 5230 4208
rect 13817 4199 13875 4205
rect 13817 4165 13829 4199
rect 13863 4196 13875 4199
rect 14185 4199 14243 4205
rect 14185 4196 14197 4199
rect 13863 4168 14197 4196
rect 13863 4165 13875 4168
rect 13817 4159 13875 4165
rect 14185 4165 14197 4168
rect 14231 4165 14243 4199
rect 14185 4159 14243 4165
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2222 3924 2228 3936
rect 1903 3896 2228 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2222 3884 2228 3896
rect 2280 3924 2286 3936
rect 3344 3924 3372 4091
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5307 4100 6914 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3752 4032 3985 4060
rect 3752 4020 3758 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 4246 4020 4252 4072
rect 4304 4020 4310 4072
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 4264 3992 4292 4020
rect 3559 3964 4292 3992
rect 4525 3995 4583 4001
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 4525 3961 4537 3995
rect 4571 3961 4583 3995
rect 6886 3992 6914 4100
rect 11790 4088 11796 4140
rect 11848 4088 11854 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 11900 4100 12909 4128
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11900 4060 11928 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 11388 4032 11928 4060
rect 11388 4020 11394 4032
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 12860 4032 13492 4060
rect 12860 4020 12866 4032
rect 12342 3992 12348 4004
rect 6886 3964 12348 3992
rect 4525 3955 4583 3961
rect 2280 3896 3372 3924
rect 2280 3884 2286 3896
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4540 3924 4568 3955
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 13464 3992 13492 4032
rect 13538 4020 13544 4072
rect 13596 4020 13602 4072
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 14108 3992 14136 4091
rect 13464 3964 14136 3992
rect 4304 3896 4568 3924
rect 4304 3884 4310 3896
rect 11882 3884 11888 3936
rect 11940 3884 11946 3936
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13262 3924 13268 3936
rect 13127 3896 13268 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 934 3680 940 3732
rect 992 3720 998 3732
rect 1489 3723 1547 3729
rect 1489 3720 1501 3723
rect 992 3692 1501 3720
rect 992 3680 998 3692
rect 1489 3689 1501 3692
rect 1535 3689 1547 3723
rect 1489 3683 1547 3689
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 11790 3720 11796 3732
rect 2004 3692 11796 3720
rect 2004 3680 2010 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12802 3680 12808 3732
rect 12860 3680 12866 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14415 3692 14872 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14844 3664 14872 3692
rect 11330 3612 11336 3664
rect 11388 3612 11394 3664
rect 14826 3612 14832 3664
rect 14884 3612 14890 3664
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2961 3587 3019 3593
rect 2961 3584 2973 3587
rect 2280 3556 2973 3584
rect 2280 3544 2286 3556
rect 2961 3553 2973 3556
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 11164 3556 11560 3584
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 1636 3488 2053 3516
rect 1636 3476 1642 3488
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2556 3488 2697 3516
rect 2556 3476 2562 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 11164 3525 11192 3556
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11532 3516 11560 3556
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13872 3556 13921 3584
rect 13872 3544 13878 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 12802 3516 12808 3528
rect 11532 3488 12808 3516
rect 11425 3479 11483 3485
rect 1762 3408 1768 3460
rect 1820 3408 1826 3460
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 4246 3448 4252 3460
rect 2004 3420 4252 3448
rect 2004 3408 2010 3420
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 4801 3451 4859 3457
rect 4801 3417 4813 3451
rect 4847 3417 4859 3451
rect 4801 3411 4859 3417
rect 4893 3451 4951 3457
rect 4893 3417 4905 3451
rect 4939 3448 4951 3451
rect 5077 3451 5135 3457
rect 5077 3448 5089 3451
rect 4939 3420 5089 3448
rect 4939 3417 4951 3420
rect 4893 3411 4951 3417
rect 5077 3417 5089 3420
rect 5123 3417 5135 3451
rect 11440 3448 11468 3479
rect 12802 3476 12808 3488
rect 12860 3516 12866 3528
rect 13446 3516 13452 3528
rect 12860 3488 13452 3516
rect 12860 3476 12866 3488
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 5077 3411 5135 3417
rect 11164 3420 11468 3448
rect 11692 3451 11750 3457
rect 1118 3340 1124 3392
rect 1176 3380 1182 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 1176 3352 2145 3380
rect 1176 3340 1182 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 3602 3340 3608 3392
rect 3660 3340 3666 3392
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4816 3380 4844 3411
rect 11164 3392 11192 3420
rect 11692 3417 11704 3451
rect 11738 3448 11750 3451
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 11738 3420 12909 3448
rect 11738 3417 11750 3420
rect 11692 3411 11750 3417
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 12897 3411 12955 3417
rect 4203 3352 4844 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 11146 3340 11152 3392
rect 11204 3340 11210 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 14200 3380 14228 3479
rect 11664 3352 14228 3380
rect 11664 3340 11670 3352
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1820 3148 1869 3176
rect 1820 3136 1826 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 1857 3139 1915 3145
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 2406 3176 2412 3188
rect 2271 3148 2412 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 2498 3136 2504 3188
rect 2556 3136 2562 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3234 3176 3240 3188
rect 3099 3148 3240 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4028 3148 4445 3176
rect 4028 3136 4034 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 4706 3136 4712 3188
rect 4764 3136 4770 3188
rect 11606 3136 11612 3188
rect 11664 3136 11670 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 11940 3148 12572 3176
rect 11940 3136 11946 3148
rect 2516 3108 2544 3136
rect 2056 3080 2544 3108
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2056 3049 2084 3080
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2280 3012 2329 3040
rect 2280 3000 2286 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 3804 3040 3832 3136
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 7650 3108 7656 3120
rect 4387 3080 7656 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 7650 3068 7656 3080
rect 7708 3108 7714 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7708 3080 7849 3108
rect 7708 3068 7714 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 3804 3012 4629 3040
rect 2317 3003 2375 3009
rect 4617 3009 4629 3012
rect 4663 3040 4675 3043
rect 4798 3040 4804 3052
rect 4663 3012 4804 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 11146 3040 11152 3052
rect 9631 3012 11152 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 11146 3000 11152 3012
rect 11204 3040 11210 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11204 3012 11529 3040
rect 11204 3000 11210 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 4816 2972 4844 3000
rect 11624 2972 11652 3136
rect 11784 3111 11842 3117
rect 11784 3077 11796 3111
rect 11830 3108 11842 3111
rect 12434 3108 12440 3120
rect 11830 3080 12440 3108
rect 11830 3077 11842 3080
rect 11784 3071 11842 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12544 3040 12572 3148
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12860 3148 12909 3176
rect 12860 3136 12866 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 12897 3139 12955 3145
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12544 3012 13001 3040
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13280 3040 13308 3136
rect 13219 3012 13308 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 4816 2944 11652 2972
rect 13722 2932 13728 2984
rect 13780 2932 13786 2984
rect 13906 2932 13912 2984
rect 13964 2932 13970 2984
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 3142 2904 3148 2916
rect 1627 2876 3148 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 5626 2904 5632 2916
rect 3476 2876 5632 2904
rect 3476 2864 3482 2876
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 13630 2864 13636 2916
rect 13688 2904 13694 2916
rect 14093 2907 14151 2913
rect 14093 2904 14105 2907
rect 13688 2876 14105 2904
rect 13688 2864 13694 2876
rect 14093 2873 14105 2876
rect 14139 2873 14151 2907
rect 14093 2867 14151 2873
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 3050 2836 3056 2848
rect 2455 2808 3056 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 15010 2836 15016 2848
rect 13320 2808 15016 2836
rect 13320 2796 13326 2808
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 1670 2592 1676 2644
rect 1728 2592 1734 2644
rect 2038 2592 2044 2644
rect 2096 2592 2102 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3694 2632 3700 2644
rect 3559 2604 3700 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 4798 2592 4804 2644
rect 4856 2592 4862 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 4948 2604 5273 2632
rect 4948 2592 4954 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5776 2604 6377 2632
rect 5776 2592 5782 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7064 2604 7389 2632
rect 7064 2592 7070 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8352 2604 8953 2632
rect 8352 2592 8358 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9950 2592 9956 2644
rect 10008 2592 10014 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11112 2604 11529 2632
rect 11112 2592 11118 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 12492 2604 12909 2632
rect 12492 2592 12498 2604
rect 12897 2601 12909 2604
rect 12943 2601 12955 2635
rect 12897 2595 12955 2601
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 13722 2632 13728 2644
rect 13587 2604 13728 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 13906 2632 13912 2644
rect 13863 2604 13912 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14182 2592 14188 2644
rect 14240 2592 14246 2644
rect 1688 2564 1716 2592
rect 2317 2567 2375 2573
rect 2317 2564 2329 2567
rect 1688 2536 2329 2564
rect 2317 2533 2329 2536
rect 2363 2533 2375 2567
rect 4816 2564 4844 2592
rect 5169 2567 5227 2573
rect 5169 2564 5181 2567
rect 4816 2536 5181 2564
rect 2317 2527 2375 2533
rect 5169 2533 5181 2536
rect 5215 2533 5227 2567
rect 5169 2527 5227 2533
rect 12529 2567 12587 2573
rect 12529 2533 12541 2567
rect 12575 2533 12587 2567
rect 12529 2527 12587 2533
rect 2240 2468 2636 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1854 2428 1860 2440
rect 1719 2400 1860 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2240 2437 2268 2468
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2130 2320 2136 2372
rect 2188 2360 2194 2372
rect 2516 2360 2544 2391
rect 2188 2332 2544 2360
rect 2608 2360 2636 2468
rect 3050 2456 3056 2508
rect 3108 2456 3114 2508
rect 3142 2456 3148 2508
rect 3200 2456 3206 2508
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3292 2468 3801 2496
rect 3292 2456 3298 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12544 2496 12572 2527
rect 14182 2496 14188 2508
rect 12400 2468 12572 2496
rect 13096 2468 14188 2496
rect 12400 2456 12406 2468
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3160 2428 3188 2456
rect 2915 2400 3188 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4045 2431 4103 2437
rect 4045 2428 4057 2431
rect 3660 2400 4057 2428
rect 3660 2388 3666 2400
rect 4045 2397 4057 2400
rect 4091 2397 4103 2431
rect 4045 2391 4103 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 4948 2400 5457 2428
rect 4948 2388 4954 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6052 2400 6561 2428
rect 6052 2388 6058 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7340 2400 7573 2428
rect 7340 2388 7346 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8628 2400 9137 2428
rect 8628 2388 8634 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9916 2400 10149 2428
rect 9916 2388 9922 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11204 2400 11713 2428
rect 11204 2388 11210 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12268 2360 12296 2391
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 13096 2437 13124 2468
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12492 2400 12725 2428
rect 12492 2388 12498 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13170 2388 13176 2440
rect 13228 2388 13234 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13372 2400 13461 2428
rect 13262 2360 13268 2372
rect 2608 2332 5580 2360
rect 12268 2332 13268 2360
rect 2188 2320 2194 2332
rect 5552 2301 5580 2332
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 12710 2292 12716 2304
rect 12483 2264 12716 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 13372 2301 13400 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13717 2433 13775 2439
rect 13717 2430 13729 2433
rect 13449 2391 13507 2397
rect 13556 2402 13729 2430
rect 13556 2360 13584 2402
rect 13717 2399 13729 2402
rect 13763 2399 13775 2433
rect 13717 2393 13775 2399
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 13464 2332 13584 2360
rect 13464 2304 13492 2332
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13446 2252 13452 2304
rect 13504 2252 13510 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14108 2292 14136 2391
rect 13596 2264 14136 2292
rect 13596 2252 13602 2264
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
<< via1 >>
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 13728 17323 13780 17332
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 1032 17212 1084 17264
rect 940 17144 992 17196
rect 2780 17144 2832 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1860 16983 1912 16992
rect 1860 16949 1869 16983
rect 1869 16949 1903 16983
rect 1903 16949 1912 16983
rect 1860 16940 1912 16949
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 1584 16736 1636 16788
rect 940 16532 992 16584
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 14372 16532 14424 16584
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 1032 15376 1084 15428
rect 14188 15376 14240 15428
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 940 14968 992 15020
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 1768 14764 1820 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 13728 13812 13780 13864
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 14832 13404 14884 13456
rect 1032 13336 1084 13388
rect 1860 13268 1912 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 1860 12384 1912 12436
rect 1768 12180 1820 12232
rect 1676 12044 1728 12096
rect 14188 12044 14240 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 940 11704 992 11756
rect 1032 11636 1084 11688
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 13820 10752 13872 10804
rect 940 10616 992 10668
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 14832 10140 14884 10192
rect 13912 10004 13964 10056
rect 10600 9936 10652 9988
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 10600 9163 10652 9172
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 11060 8916 11112 8968
rect 940 8848 992 8900
rect 1768 8891 1820 8900
rect 1768 8857 1777 8891
rect 1777 8857 1811 8891
rect 1811 8857 1820 8891
rect 1768 8848 1820 8857
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 1768 8576 1820 8628
rect 1676 8508 1728 8560
rect 5540 8440 5592 8492
rect 9956 8440 10008 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 14464 8304 14516 8356
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 5540 7488 5592 7540
rect 6828 7352 6880 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 940 7148 992 7200
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 1584 6808 1636 6860
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 14372 6740 14424 6792
rect 940 6672 992 6724
rect 5540 6672 5592 6724
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 13912 6647 13964 6656
rect 13912 6613 13921 6647
rect 13921 6613 13955 6647
rect 13955 6613 13964 6647
rect 13912 6604 13964 6613
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 2044 6400 2096 6452
rect 11704 6400 11756 6452
rect 13452 6400 13504 6452
rect 14188 6400 14240 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 13268 6332 13320 6384
rect 13912 6332 13964 6384
rect 13084 6264 13136 6316
rect 12808 6196 12860 6248
rect 14188 6128 14240 6180
rect 3424 6060 3476 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 1676 5856 1728 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 11796 5856 11848 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13268 5856 13320 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 4712 5788 4764 5840
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 5540 5720 5592 5772
rect 3148 5584 3200 5636
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 12624 5788 12676 5840
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 3792 5516 3844 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 13636 5652 13688 5704
rect 13820 5584 13872 5636
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 11796 5312 11848 5364
rect 12440 5312 12492 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 2412 5287 2464 5296
rect 2412 5253 2421 5287
rect 2421 5253 2455 5287
rect 2455 5253 2464 5287
rect 2412 5244 2464 5253
rect 2044 5176 2096 5228
rect 3148 5176 3200 5228
rect 4252 5176 4304 5228
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 5540 5108 5592 5160
rect 11152 5108 11204 5160
rect 12716 5108 12768 5160
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 940 4972 992 5024
rect 2320 4972 2372 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 4436 4972 4488 5024
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 2504 4768 2556 4820
rect 3792 4768 3844 4820
rect 4436 4768 4488 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 3424 4632 3476 4684
rect 3792 4564 3844 4616
rect 5172 4564 5224 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 9036 4564 9088 4616
rect 1860 4496 1912 4548
rect 2320 4496 2372 4548
rect 3056 4496 3108 4548
rect 4160 4496 4212 4548
rect 12164 4496 12216 4548
rect 13544 4496 13596 4548
rect 3148 4428 3200 4480
rect 7656 4428 7708 4480
rect 12808 4428 12860 4480
rect 13820 4539 13872 4548
rect 13820 4505 13829 4539
rect 13829 4505 13863 4539
rect 13863 4505 13872 4539
rect 13820 4496 13872 4505
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 2780 4224 2832 4276
rect 3148 4156 3200 4208
rect 9036 4224 9088 4276
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 5172 4199 5224 4208
rect 5172 4165 5181 4199
rect 5181 4165 5215 4199
rect 5215 4165 5224 4199
rect 5172 4156 5224 4165
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 2228 3884 2280 3936
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 3700 4020 3752 4072
rect 4252 4020 4304 4072
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 11336 4020 11388 4072
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 4252 3884 4304 3936
rect 12348 3952 12400 4004
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 13636 4020 13688 4072
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13268 3884 13320 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 940 3680 992 3732
rect 1952 3680 2004 3732
rect 11796 3680 11848 3732
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 11336 3655 11388 3664
rect 11336 3621 11345 3655
rect 11345 3621 11379 3655
rect 11379 3621 11388 3655
rect 11336 3612 11388 3621
rect 14832 3612 14884 3664
rect 2228 3544 2280 3596
rect 1584 3476 1636 3528
rect 2504 3476 2556 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 13820 3544 13872 3596
rect 1768 3451 1820 3460
rect 1768 3417 1777 3451
rect 1777 3417 1811 3451
rect 1811 3417 1820 3451
rect 1768 3408 1820 3417
rect 1952 3408 2004 3460
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 12808 3476 12860 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 1124 3340 1176 3392
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 11152 3340 11204 3392
rect 11612 3340 11664 3392
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 1768 3136 1820 3188
rect 2412 3136 2464 3188
rect 2504 3136 2556 3188
rect 3240 3136 3292 3188
rect 3792 3136 3844 3188
rect 3976 3136 4028 3188
rect 4712 3179 4764 3188
rect 4712 3145 4721 3179
rect 4721 3145 4755 3179
rect 4755 3145 4764 3179
rect 4712 3136 4764 3145
rect 11612 3136 11664 3188
rect 11888 3136 11940 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2228 3000 2280 3052
rect 7656 3068 7708 3120
rect 4804 3000 4856 3052
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 11152 3000 11204 3052
rect 12440 3068 12492 3120
rect 12808 3136 12860 3188
rect 13268 3136 13320 3188
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 3148 2864 3200 2916
rect 3424 2864 3476 2916
rect 5632 2864 5684 2916
rect 13636 2907 13688 2916
rect 13636 2873 13645 2907
rect 13645 2873 13679 2907
rect 13679 2873 13688 2907
rect 13636 2864 13688 2873
rect 3056 2796 3108 2848
rect 13268 2796 13320 2848
rect 15016 2796 15068 2848
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 1676 2592 1728 2644
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 3700 2592 3752 2644
rect 4804 2592 4856 2644
rect 4896 2592 4948 2644
rect 5724 2592 5776 2644
rect 7012 2592 7064 2644
rect 8300 2592 8352 2644
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 11060 2592 11112 2644
rect 12440 2592 12492 2644
rect 13728 2592 13780 2644
rect 13912 2592 13964 2644
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 1860 2388 1912 2440
rect 2136 2320 2188 2372
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 3056 2456 3108 2465
rect 3148 2456 3200 2508
rect 3240 2456 3292 2508
rect 12348 2456 12400 2508
rect 3608 2388 3660 2440
rect 4896 2388 4948 2440
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6000 2388 6052 2440
rect 7288 2388 7340 2440
rect 8576 2388 8628 2440
rect 9864 2388 9916 2440
rect 11152 2388 11204 2440
rect 12440 2388 12492 2440
rect 14188 2456 14240 2508
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 13268 2320 13320 2372
rect 12716 2252 12768 2304
rect 13452 2252 13504 2304
rect 13544 2252 13596 2304
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
<< metal2 >>
rect 2778 18592 2834 18601
rect 2778 18527 2834 18536
rect 1030 17776 1086 17785
rect 1030 17711 1086 17720
rect 1044 17270 1072 17711
rect 1032 17264 1084 17270
rect 1032 17206 1084 17212
rect 2792 17202 2820 18527
rect 13726 18048 13782 18057
rect 13726 17983 13782 17992
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 13740 17338 13768 17983
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 952 16969 980 17138
rect 1872 17054 2084 17082
rect 1872 16998 1900 17054
rect 1584 16992 1636 16998
rect 938 16960 994 16969
rect 1584 16934 1636 16940
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 938 16895 994 16904
rect 1596 16794 1624 16934
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 940 16584 992 16590
rect 940 16526 992 16532
rect 952 16153 980 16526
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 938 16144 994 16153
rect 938 16079 994 16088
rect 1596 15502 1624 16390
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1032 15428 1084 15434
rect 1032 15370 1084 15376
rect 1044 15337 1072 15370
rect 1860 15360 1912 15366
rect 1030 15328 1086 15337
rect 1860 15302 1912 15308
rect 1030 15263 1086 15272
rect 940 15020 992 15026
rect 940 14962 992 14968
rect 952 14521 980 14962
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 938 14512 994 14521
rect 938 14447 994 14456
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1032 13388 1084 13394
rect 1032 13330 1084 13336
rect 1044 12889 1072 13330
rect 1030 12880 1086 12889
rect 1030 12815 1086 12824
rect 1780 12238 1808 14758
rect 1872 13326 1900 15302
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12442 1900 13126
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1676 12096 1728 12102
rect 938 12064 994 12073
rect 1676 12038 1728 12044
rect 938 11999 994 12008
rect 952 11762 980 11999
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 1032 11688 1084 11694
rect 1032 11630 1084 11636
rect 1044 11257 1072 11630
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1030 11248 1086 11257
rect 1030 11183 1086 11192
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10441 980 10610
rect 938 10432 994 10441
rect 938 10367 994 10376
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8809 980 8842
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 940 7200 992 7206
rect 938 7168 940 7177
rect 992 7168 994 7177
rect 938 7103 994 7112
rect 1596 6866 1624 11494
rect 1688 8566 1716 12038
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1780 8634 1808 8842
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6361 980 6666
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1688 5914 1716 6258
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 1872 5250 1900 11494
rect 1964 6798 1992 16934
rect 2056 16574 2084 17054
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12944 16827 13252 16836
rect 2056 16546 2176 16574
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6458 2084 6598
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2148 6338 2176 16546
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 13740 13326 13768 13806
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 13832 10810 13860 17138
rect 14372 16584 14424 16590
rect 14370 16552 14372 16561
rect 14424 16552 14426 16561
rect 14370 16487 14426 16496
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14200 15026 14228 15370
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14372 14816 14424 14822
rect 14370 14784 14372 14793
rect 14424 14784 14426 14793
rect 14370 14719 14426 14728
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14844 13297 14872 13398
rect 14830 13288 14886 13297
rect 14830 13223 14886 13232
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13924 10062 13952 13126
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11762 14228 12038
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14372 11552 14424 11558
rect 14370 11520 14372 11529
rect 14424 11520 14426 11529
rect 14370 11455 14426 11464
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 13912 10056 13964 10062
rect 14844 10033 14872 10134
rect 13912 9998 13964 10004
rect 14830 10024 14886 10033
rect 10600 9988 10652 9994
rect 14830 9959 14886 9968
rect 10600 9930 10652 9936
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 10612 9178 10640 9930
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 5552 7546 5580 8434
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6840 7002 6868 7346
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 2056 6310 2176 6338
rect 2056 5710 2084 6310
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 2412 5296 2464 5302
rect 1872 5222 1992 5250
rect 2412 5238 2464 5244
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4729 980 4966
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 938 3904 994 3913
rect 938 3839 994 3848
rect 952 3738 980 3839
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1124 3392 1176 3398
rect 1124 3334 1176 3340
rect 1136 3097 1164 3334
rect 1122 3088 1178 3097
rect 1122 3023 1178 3032
rect 1596 2650 1624 3470
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 3194 1808 3402
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 2650 1716 2994
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1872 2446 1900 4490
rect 1964 3738 1992 5222
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1964 3058 1992 3402
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2056 2650 2084 5170
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4554 2360 4966
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3602 2268 3878
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3058 2268 3538
rect 2424 3194 2452 5238
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2516 3534 2544 4762
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4282 2820 4626
rect 3068 4554 3096 5510
rect 3160 5234 3188 5578
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3436 4690 3464 6054
rect 5552 5914 5580 6666
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 3160 4214 3188 4422
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 3194 2544 3334
rect 3252 3194 3280 4082
rect 3712 4078 3740 4966
rect 3804 4826 3832 5510
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3804 4622 3832 4762
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 3068 2514 3096 2790
rect 3160 2514 3188 2858
rect 3252 2514 3280 3130
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2136 2372 2188 2378
rect 2136 2314 2188 2320
rect 2148 800 2176 2314
rect 3436 800 3464 2858
rect 3620 2446 3648 3334
rect 3712 2650 3740 4014
rect 3804 3194 3832 4082
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3194 4016 3470
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 4066 2272 4122 2281
rect 4172 2258 4200 4490
rect 4264 4078 4292 5170
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4826 4476 4966
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 3466 4292 3878
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 4724 3194 4752 5782
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5166 5580 5714
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4622 5580 5102
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5184 4214 5212 4558
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4816 2650 4844 2994
rect 4908 2650 4936 2994
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4896 2440 4948 2446
rect 4122 2230 4200 2258
rect 4724 2400 4896 2428
rect 4066 2207 4122 2216
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 4724 800 4752 2400
rect 5644 2428 5672 2858
rect 5736 2650 5764 5646
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 6090 2683 6398 2692
rect 7024 2650 7052 6734
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 3126 7696 4422
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 8312 2650 8340 7346
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9048 4282 9076 4558
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 9968 2650 9996 8434
rect 11072 2650 11100 8910
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 8265 14504 8298
rect 14462 8256 14518 8265
rect 12944 8188 13252 8197
rect 14462 8191 14518 8200
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 14188 6792 14240 6798
rect 14372 6792 14424 6798
rect 14188 6734 14240 6740
rect 14370 6760 14372 6769
rect 14424 6760 14426 6769
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11716 6458 11744 6598
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 13280 6390 13308 6734
rect 13464 6458 13492 6734
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13924 6390 13952 6598
rect 14200 6458 14228 6734
rect 14370 6695 14426 6704
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 11808 5914 11836 6258
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 13096 6202 13124 6258
rect 12820 5914 12848 6190
rect 13096 6174 13308 6202
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 13280 5914 13308 6174
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14200 5914 14228 6122
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11808 5370 11836 5510
rect 12452 5370 12480 5646
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11164 3398 11192 5102
rect 12636 4826 12664 5782
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13648 5234 13676 5646
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5370 13860 5578
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 12176 4282 12204 4490
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3670 11376 4014
rect 11808 3738 11836 4082
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11164 3058 11192 3334
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 11624 3194 11652 3334
rect 11900 3194 11928 3878
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 12360 2514 12388 3946
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12452 2650 12480 3062
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 5724 2440 5776 2446
rect 5644 2400 5724 2428
rect 4896 2382 4948 2388
rect 5724 2382 5776 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 6012 800 6040 2382
rect 7300 800 7328 2382
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 8588 800 8616 2382
rect 9876 800 9904 2382
rect 11164 800 11192 2382
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 12452 800 12480 2382
rect 12728 2310 12756 5102
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4078 12848 4422
rect 13556 4078 13584 4490
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 12820 3738 12848 4014
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12820 3194 12848 3470
rect 13280 3194 13308 3878
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 13280 2530 13308 2790
rect 13188 2502 13308 2530
rect 13188 2446 13216 2502
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 2134 0 2190 800
rect 3422 0 3478 800
rect 4710 0 4766 800
rect 5998 0 6054 800
rect 7286 0 7342 800
rect 8574 0 8630 800
rect 9862 0 9918 800
rect 11150 0 11206 800
rect 12438 0 12494 800
rect 13280 762 13308 2314
rect 13464 2310 13492 3470
rect 13556 2310 13584 4014
rect 13648 2922 13676 4014
rect 13832 3602 13860 4490
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13740 2650 13768 2926
rect 13924 2650 13952 2926
rect 14200 2650 14228 5170
rect 14372 5024 14424 5030
rect 14370 4992 14372 5001
rect 14424 4992 14426 5001
rect 14370 4927 14426 4936
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 3505 14872 3606
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14200 1737 14228 2450
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 14186 1728 14242 1737
rect 14186 1663 14242 1672
rect 13648 870 13768 898
rect 13648 762 13676 870
rect 13740 800 13768 870
rect 15028 800 15056 2790
rect 13280 734 13676 762
rect 13726 0 13782 800
rect 15014 0 15070 800
<< via2 >>
rect 2778 18536 2834 18592
rect 1030 17720 1086 17776
rect 13726 17992 13782 18048
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 938 16904 994 16960
rect 938 16088 994 16144
rect 1030 15272 1086 15328
rect 938 14456 994 14512
rect 1398 13640 1454 13696
rect 1030 12824 1086 12880
rect 938 12008 994 12064
rect 1030 11192 1086 11248
rect 938 10376 994 10432
rect 1490 9560 1546 9616
rect 938 8744 994 8800
rect 1490 8200 1546 8256
rect 938 7148 940 7168
rect 940 7148 992 7168
rect 992 7148 994 7168
rect 938 7112 994 7148
rect 938 6296 994 6352
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 14370 16532 14372 16552
rect 14372 16532 14424 16552
rect 14424 16532 14426 16552
rect 14370 16496 14426 16532
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14370 14764 14372 14784
rect 14372 14764 14424 14784
rect 14424 14764 14426 14784
rect 14370 14728 14426 14764
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14830 13232 14886 13288
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14370 11500 14372 11520
rect 14372 11500 14424 11520
rect 14424 11500 14426 11520
rect 14370 11464 14426 11500
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14830 9968 14886 10024
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 938 4664 994 4720
rect 938 3848 994 3904
rect 1122 3032 1178 3088
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4066 2216 4122 2272
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14462 8200 14518 8256
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 14370 6740 14372 6760
rect 14372 6740 14424 6760
rect 14424 6740 14426 6760
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 14370 6704 14426 6740
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14370 4972 14372 4992
rect 14372 4972 14424 4992
rect 14424 4972 14426 4992
rect 14370 4936 14426 4972
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14830 3440 14886 3496
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 14186 1672 14242 1728
<< metal3 >>
rect 0 18594 800 18624
rect 2773 18594 2839 18597
rect 0 18592 2839 18594
rect 0 18536 2778 18592
rect 2834 18536 2839 18592
rect 0 18534 2839 18536
rect 0 18504 800 18534
rect 2773 18531 2839 18534
rect 13721 18050 13787 18053
rect 15200 18050 16000 18080
rect 13721 18048 16000 18050
rect 13721 17992 13726 18048
rect 13782 17992 16000 18048
rect 13721 17990 16000 17992
rect 13721 17987 13787 17990
rect 15200 17960 16000 17990
rect 0 17778 800 17808
rect 1025 17778 1091 17781
rect 0 17776 1091 17778
rect 0 17720 1030 17776
rect 1086 17720 1091 17776
rect 0 17718 1091 17720
rect 0 17688 800 17718
rect 1025 17715 1091 17718
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 14653 17375 14969 17376
rect 0 16962 800 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 800 16902
rect 933 16899 999 16902
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 12940 16831 13256 16832
rect 14365 16554 14431 16557
rect 14365 16552 15210 16554
rect 14365 16496 14370 16552
rect 14426 16496 15210 16552
rect 14365 16494 15210 16496
rect 14365 16491 14431 16494
rect 15150 16448 15210 16494
rect 15150 16358 16000 16448
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 15200 16328 16000 16358
rect 14653 16287 14969 16288
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 12940 15743 13256 15744
rect 0 15330 800 15360
rect 1025 15330 1091 15333
rect 0 15328 1091 15330
rect 0 15272 1030 15328
rect 1086 15272 1091 15328
rect 0 15270 1091 15272
rect 0 15240 800 15270
rect 1025 15267 1091 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 14653 15199 14969 15200
rect 14365 14786 14431 14789
rect 15200 14786 16000 14816
rect 14365 14784 16000 14786
rect 14365 14728 14370 14784
rect 14426 14728 16000 14784
rect 14365 14726 16000 14728
rect 14365 14723 14431 14726
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 15200 14696 16000 14726
rect 12940 14655 13256 14656
rect 0 14514 800 14544
rect 933 14514 999 14517
rect 0 14512 999 14514
rect 0 14456 938 14512
rect 994 14456 999 14512
rect 0 14454 999 14456
rect 0 14424 800 14454
rect 933 14451 999 14454
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 14653 14111 14969 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 14825 13290 14891 13293
rect 14825 13288 15210 13290
rect 14825 13232 14830 13288
rect 14886 13232 15210 13288
rect 14825 13230 15210 13232
rect 14825 13227 14891 13230
rect 15150 13184 15210 13230
rect 15150 13094 16000 13184
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 15200 13064 16000 13094
rect 14653 13023 14969 13024
rect 0 12882 800 12912
rect 1025 12882 1091 12885
rect 0 12880 1091 12882
rect 0 12824 1030 12880
rect 1086 12824 1091 12880
rect 0 12822 1091 12824
rect 0 12792 800 12822
rect 1025 12819 1091 12822
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 12940 12479 13256 12480
rect 0 12066 800 12096
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 0 11976 800 12006
rect 933 12003 999 12006
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 14653 11935 14969 11936
rect 14365 11522 14431 11525
rect 15200 11522 16000 11552
rect 14365 11520 16000 11522
rect 14365 11464 14370 11520
rect 14426 11464 16000 11520
rect 14365 11462 16000 11464
rect 14365 11459 14431 11462
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 15200 11432 16000 11462
rect 12940 11391 13256 11392
rect 0 11250 800 11280
rect 1025 11250 1091 11253
rect 0 11248 1091 11250
rect 0 11192 1030 11248
rect 1086 11192 1091 11248
rect 0 11190 1091 11192
rect 0 11160 800 11190
rect 1025 11187 1091 11190
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 14653 10847 14969 10848
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 12940 10303 13256 10304
rect 14825 10026 14891 10029
rect 14825 10024 15210 10026
rect 14825 9968 14830 10024
rect 14886 9968 15210 10024
rect 14825 9966 15210 9968
rect 14825 9963 14891 9966
rect 15150 9920 15210 9966
rect 15150 9830 16000 9920
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 15200 9800 16000 9830
rect 14653 9759 14969 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 12940 9215 13256 9216
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 14653 8671 14969 8672
rect 1485 8258 1551 8261
rect 798 8256 1551 8258
rect 798 8200 1490 8256
rect 1546 8200 1551 8256
rect 798 8198 1551 8200
rect 798 8016 858 8198
rect 1485 8195 1551 8198
rect 14457 8258 14523 8261
rect 15200 8258 16000 8288
rect 14457 8256 16000 8258
rect 14457 8200 14462 8256
rect 14518 8200 16000 8256
rect 14457 8198 16000 8200
rect 14457 8195 14523 8198
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 15200 8168 16000 8198
rect 12940 8127 13256 8128
rect 0 7926 858 8016
rect 0 7896 800 7926
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 14653 7583 14969 7584
rect 0 7170 800 7200
rect 933 7170 999 7173
rect 0 7168 999 7170
rect 0 7112 938 7168
rect 994 7112 999 7168
rect 0 7110 999 7112
rect 0 7080 800 7110
rect 933 7107 999 7110
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 12940 7039 13256 7040
rect 14365 6762 14431 6765
rect 14365 6760 15210 6762
rect 14365 6704 14370 6760
rect 14426 6704 15210 6760
rect 14365 6702 15210 6704
rect 14365 6699 14431 6702
rect 15150 6656 15210 6702
rect 15150 6566 16000 6656
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 15200 6536 16000 6566
rect 14653 6495 14969 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 14653 5407 14969 5408
rect 14365 4994 14431 4997
rect 15200 4994 16000 5024
rect 14365 4992 16000 4994
rect 14365 4936 14370 4992
rect 14426 4936 16000 4992
rect 14365 4934 16000 4936
rect 14365 4931 14431 4934
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 15200 4904 16000 4934
rect 12940 4863 13256 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 14825 3498 14891 3501
rect 14825 3496 15210 3498
rect 14825 3440 14830 3496
rect 14886 3440 15210 3496
rect 14825 3438 15210 3440
rect 14825 3435 14891 3438
rect 15150 3392 15210 3438
rect 15150 3302 16000 3392
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 15200 3272 16000 3302
rect 14653 3231 14969 3232
rect 0 3090 800 3120
rect 1117 3090 1183 3093
rect 0 3088 1183 3090
rect 0 3032 1122 3088
rect 1178 3032 1183 3088
rect 0 3030 1183 3032
rect 0 3000 800 3030
rect 1117 3027 1183 3030
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 0 2274 800 2304
rect 4061 2274 4127 2277
rect 0 2272 4127 2274
rect 0 2216 4066 2272
rect 4122 2216 4127 2272
rect 0 2214 4127 2216
rect 0 2184 800 2214
rect 4061 2211 4127 2214
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 14181 1730 14247 1733
rect 15200 1730 16000 1760
rect 14181 1728 16000 1730
rect 14181 1672 14186 1728
rect 14242 1672 16000 1728
rect 14181 1670 16000 1672
rect 14181 1667 14247 1670
rect 15200 1640 16000 1670
<< via3 >>
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
<< metal4 >>
rect 2657 16896 2977 17456
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 2128 2977 2688
rect 4370 17440 4690 17456
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 2128 4690 2144
rect 6084 16896 6404 17456
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 6084 2128 6404 2688
rect 7797 17440 8117 17456
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 2128 8117 2144
rect 9511 16896 9831 17456
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 2128 9831 2688
rect 11224 17440 11544 17456
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 2128 11544 2144
rect 12938 16896 13258 17456
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12938 15808 13258 16832
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12938 8192 13258 9216
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 2128 13258 2688
rect 14651 17440 14971 17456
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 2128 14971 2144
use sky130_fd_sc_hd__inv_2  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp 1688980957
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 1688980957
transform -1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform -1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _039_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform -1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform -1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform -1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform -1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform -1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform -1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp 1688980957
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _054_
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1688980957
transform 1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1688980957
transform -1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1688980957
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1688980957
transform -1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1688980957
transform -1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1688980957
transform -1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _064_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _065_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _066_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _067_
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _068_
timestamp 1688980957
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _069_
timestamp 1688980957
transform -1 0 10948 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _070_
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _071_
timestamp 1688980957
transform -1 0 3312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform -1 0 13984 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp 1688980957
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp 1688980957
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp 1688980957
transform 1 0 1564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _090_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _091_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14076 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _092_
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _093_
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _093__43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _094_
timestamp 1688980957
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _094__44
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _095_
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _096_
timestamp 1688980957
transform -1 0 13432 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _097_
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _098__45
timestamp 1688980957
transform -1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _098_
timestamp 1688980957
transform 1 0 2208 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _099_
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _100_
timestamp 1688980957
transform -1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _101_
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _102_
timestamp 1688980957
transform 1 0 3220 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _103__46
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _103_
timestamp 1688980957
transform -1 0 5060 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _104_
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _105_
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk
timestamp 1688980957
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_16
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_71 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_88
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_116
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_120
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_144 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_42
timestamp 1688980957
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_145
timestamp 1688980957
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_18
timestamp 1688980957
transform 1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_46
timestamp 1688980957
transform 1 0 5336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_70
timestamp 1688980957
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_46
timestamp 1688980957
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1688980957
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_131
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_144
timestamp 1688980957
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_49
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_57
timestamp 1688980957
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_126
timestamp 1688980957
transform 1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_144
timestamp 1688980957
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_21
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_34
timestamp 1688980957
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_46
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_65
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_89
timestamp 1688980957
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1688980957
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_16
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_23
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 1688980957
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_63
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_75
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_124
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_17
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_41
timestamp 1688980957
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_127
timestamp 1688980957
transform 1 0 12788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_12
timestamp 1688980957
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_24
timestamp 1688980957
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_61
timestamp 1688980957
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_113
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_117
timestamp 1688980957
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_129
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_33
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_75
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_79
timestamp 1688980957
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_91
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_103
timestamp 1688980957
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_145
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_106
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_118
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_130
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_9
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_21
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1688980957
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_143
timestamp 1688980957
transform 1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_145
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1688980957
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_141
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_11
timestamp 1688980957
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 1688980957
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_145
timestamp 1688980957
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 1688980957
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 1688980957
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 1688980957
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1688980957
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_145
timestamp 1688980957
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_6
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_18
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_30
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1688980957
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_11
timestamp 1688980957
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_23
timestamp 1688980957
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_145
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_145
timestamp 1688980957
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_6
timestamp 1688980957
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 1688980957
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_12
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_24
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 13616 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform -1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1688980957
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 1932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform -1 0 1932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform -1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1688980957
transform 1 0 14168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1688980957
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform -1 0 13984 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
port 0 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 1 nsew signal input
flabel metal3 s 15200 1640 16000 1760 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 15200 3272 16000 3392 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 5 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 6 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 7 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 8 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 9 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 10 nsew signal input
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 11 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 12 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 13 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 14 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 15 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 16 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 17 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 18 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 19 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 20 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 21 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 22 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 23 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 24 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 25 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 26 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 27 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 28 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 29 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 30 nsew signal input
flabel metal3 s 15200 4904 16000 5024 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 31 nsew signal tristate
flabel metal3 s 15200 6536 16000 6656 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 32 nsew signal tristate
flabel metal3 s 15200 8168 16000 8288 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 33 nsew signal tristate
flabel metal3 s 15200 9800 16000 9920 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 34 nsew signal tristate
flabel metal3 s 15200 11432 16000 11552 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 35 nsew signal tristate
flabel metal3 s 15200 13064 16000 13184 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 36 nsew signal tristate
flabel metal3 s 15200 14696 16000 14816 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 37 nsew signal tristate
flabel metal3 s 15200 16328 16000 16448 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 38 nsew signal tristate
flabel metal3 s 15200 17960 16000 18080 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 39 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 40 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 41 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 prog_clk
port 42 nsew signal input
flabel metal4 s 2657 2128 2977 17456 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 6084 2128 6404 17456 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 9511 2128 9831 17456 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 12938 2128 13258 17456 0 FreeSans 1920 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 4370 2128 4690 17456 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 7797 2128 8117 17456 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 11224 2128 11544 17456 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 14651 2128 14971 17456 0 FreeSans 1920 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 7958 16864 7958 16864 0 vdd
rlabel via1 8037 17408 8037 17408 0 vss
rlabel metal1 4232 3162 4232 3162 0 _000_
rlabel metal1 3910 3978 3910 3978 0 _001_
rlabel metal1 2024 5882 2024 5882 0 _002_
rlabel metal1 2070 3060 2070 3060 0 _003_
rlabel metal1 11776 5882 11776 5882 0 _004_
rlabel metal1 13524 5882 13524 5882 0 _005_
rlabel metal1 14306 4624 14306 4624 0 _006_
rlabel metal2 11362 3842 11362 3842 0 _007_
rlabel metal1 13892 2618 13892 2618 0 _008_
rlabel metal1 14030 4182 14030 4182 0 _009_
rlabel metal1 13248 3026 13248 3026 0 _010_
rlabel metal1 13754 4488 13754 4488 0 _011_
rlabel metal1 13294 6426 13294 6426 0 _012_
rlabel metal1 12282 6188 12282 6188 0 _013_
rlabel metal1 13386 5746 13386 5746 0 _014_
rlabel metal2 14214 6018 14214 6018 0 _015_
rlabel metal1 2346 3162 2346 3162 0 _016_
rlabel metal1 2024 6222 2024 6222 0 _017_
rlabel metal1 5290 4658 5290 4658 0 _018_
rlabel metal1 3266 4522 3266 4522 0 _019_
rlabel metal1 3450 5100 3450 5100 0 _020_
rlabel metal1 4830 3400 4830 3400 0 _021_
rlabel metal1 3910 4182 3910 4182 0 _022_
rlabel metal2 3082 2652 3082 2652 0 _023_
rlabel metal2 13754 823 13754 823 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 15042 1792 15042 1792 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 13110 2448 13110 2448 0 ccff_head
rlabel metal1 14628 3706 14628 3706 0 ccff_tail
rlabel metal3 820 10404 820 10404 0 chanx_left_in[0]
rlabel metal3 866 11220 866 11220 0 chanx_left_in[1]
rlabel metal3 820 12036 820 12036 0 chanx_left_in[2]
rlabel metal3 866 12852 866 12852 0 chanx_left_in[3]
rlabel metal3 1050 13668 1050 13668 0 chanx_left_in[4]
rlabel metal3 820 14484 820 14484 0 chanx_left_in[5]
rlabel metal3 866 15300 866 15300 0 chanx_left_in[6]
rlabel metal3 820 16116 820 16116 0 chanx_left_in[7]
rlabel metal3 820 16932 820 16932 0 chanx_left_in[8]
rlabel metal3 912 3060 912 3060 0 chanx_left_out[0]
rlabel metal3 820 3876 820 3876 0 chanx_left_out[1]
rlabel metal3 820 4692 820 4692 0 chanx_left_out[2]
rlabel metal3 1096 5508 1096 5508 0 chanx_left_out[3]
rlabel metal3 820 6324 820 6324 0 chanx_left_out[4]
rlabel metal3 820 7140 820 7140 0 chanx_left_out[5]
rlabel metal3 751 7956 751 7956 0 chanx_left_out[6]
rlabel metal3 820 8772 820 8772 0 chanx_left_out[7]
rlabel metal3 1096 9588 1096 9588 0 chanx_left_out[8]
rlabel metal2 2162 1554 2162 1554 0 chany_bottom_in[0]
rlabel metal2 3450 1826 3450 1826 0 chany_bottom_in[1]
rlabel metal2 4738 1588 4738 1588 0 chany_bottom_in[2]
rlabel metal2 6026 1588 6026 1588 0 chany_bottom_in[3]
rlabel metal2 7314 1588 7314 1588 0 chany_bottom_in[4]
rlabel metal2 8602 1588 8602 1588 0 chany_bottom_in[5]
rlabel metal2 9890 1588 9890 1588 0 chany_bottom_in[6]
rlabel metal2 11178 1588 11178 1588 0 chany_bottom_in[7]
rlabel metal2 12466 1588 12466 1588 0 chany_bottom_in[8]
rlabel via2 14398 4981 14398 4981 0 chany_bottom_out[0]
rlabel via2 14398 6749 14398 6749 0 chany_bottom_out[1]
rlabel metal1 14444 8330 14444 8330 0 chany_bottom_out[2]
rlabel metal1 14628 10234 14628 10234 0 chany_bottom_out[3]
rlabel via2 14398 11509 14398 11509 0 chany_bottom_out[4]
rlabel metal1 14628 13498 14628 13498 0 chany_bottom_out[5]
rlabel via2 14398 14773 14398 14773 0 chany_bottom_out[6]
rlabel via2 14398 16541 14398 16541 0 chany_bottom_out[7]
rlabel metal2 13754 17663 13754 17663 0 chany_bottom_out[8]
rlabel metal1 7774 3094 7774 3094 0 clknet_0_prog_clk
rlabel metal1 3266 4182 3266 4182 0 clknet_1_0__leaf_prog_clk
rlabel metal1 10580 3026 10580 3026 0 clknet_1_1__leaf_prog_clk
rlabel metal3 866 17748 866 17748 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1740 18564 1740 18564 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 12880 3162 12880 3162 0 mem_bottom_track_1.DFF_0_.Q
rlabel metal1 13156 4046 13156 4046 0 mem_bottom_track_1.DFF_1_.Q
rlabel metal1 13570 5678 13570 5678 0 mem_bottom_track_3.DFF_0_.Q
rlabel metal1 12696 5338 12696 5338 0 mem_bottom_track_3.DFF_1_.Q
rlabel metal2 5566 5168 5566 5168 0 mem_left_track_1.DFF_0_.Q
rlabel metal1 3404 5678 3404 5678 0 mem_left_track_1.DFF_1_.Q
rlabel metal1 2300 3026 2300 3026 0 mem_left_track_3.DFF_0_.Q
rlabel metal1 13662 2618 13662 2618 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 12788 3026 12788 3026 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 13892 2890 13892 2890 0 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal2 13570 3162 13570 3162 0 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 13846 5474 13846 5474 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal1 12098 6324 12098 6324 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal1 12972 6222 12972 6222 0 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 14030 6290 14030 6290 0 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal2 5198 4386 5198 4386 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 2024 6290 2024 6290 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 3496 4658 3496 4658 0 mux_left_track_1.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 2392 4522 2392 4522 0 mux_left_track_1.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 3036 2414 3036 2414 0 mux_left_track_3.INVTX1_0_.out
rlabel metal1 3220 5202 3220 5202 0 mux_left_track_3.INVTX1_1_.out
rlabel metal1 3864 4046 3864 4046 0 mux_left_track_3.mux_l1_in_0_.TGATE_0_.out
rlabel metal1 3128 3434 3128 3434 0 mux_left_track_3.mux_l2_in_0_.TGATE_0_.out
rlabel metal1 12604 2278 12604 2278 0 net1
rlabel metal1 1748 13294 1748 13294 0 net10
rlabel metal2 1610 15946 1610 15946 0 net11
rlabel metal2 1610 16864 1610 16864 0 net12
rlabel metal1 2024 2550 2024 2550 0 net13
rlabel metal1 2254 2448 2254 2448 0 net14
rlabel metal1 5106 2618 5106 2618 0 net15
rlabel metal1 6072 2618 6072 2618 0 net16
rlabel metal1 7222 2618 7222 2618 0 net17
rlabel metal1 8648 2618 8648 2618 0 net18
rlabel metal1 9798 8466 9798 8466 0 net19
rlabel metal1 13432 2414 13432 2414 0 net2
rlabel metal1 11316 2618 11316 2618 0 net20
rlabel metal1 6095 4114 6095 4114 0 net21
rlabel metal2 2116 6324 2116 6324 0 net22
rlabel metal2 1978 11866 1978 11866 0 net23
rlabel metal1 4232 3026 4232 3026 0 net24
rlabel metal2 1610 3060 1610 3060 0 net25
rlabel metal1 1840 3162 1840 3162 0 net26
rlabel metal2 2070 3910 2070 3910 0 net27
rlabel metal2 4738 4488 4738 4488 0 net28
rlabel metal2 5566 6290 5566 6290 0 net29
rlabel metal1 12696 2618 12696 2618 0 net3
rlabel metal2 6854 7174 6854 7174 0 net30
rlabel metal2 5566 7990 5566 7990 0 net31
rlabel metal2 1794 8738 1794 8738 0 net32
rlabel metal2 10626 9554 10626 9554 0 net33
rlabel metal2 14214 3910 14214 3910 0 net34
rlabel metal1 14260 6426 14260 6426 0 net35
rlabel metal2 1702 10302 1702 10302 0 net36
rlabel metal1 14076 10030 14076 10030 0 net37
rlabel metal2 14214 11900 14214 11900 0 net38
rlabel metal1 1794 13192 1794 13192 0 net39
rlabel metal1 4255 10438 4255 10438 0 net4
rlabel metal1 1794 15368 1794 15368 0 net40
rlabel metal1 14076 16422 14076 16422 0 net41
rlabel metal1 13938 10778 13938 10778 0 net42
rlabel metal1 13892 3570 13892 3570 0 net43
rlabel metal1 13708 6222 13708 6222 0 net44
rlabel metal1 2254 5134 2254 5134 0 net45
rlabel metal1 5014 3434 5014 3434 0 net46
rlabel metal2 12190 4386 12190 4386 0 net47
rlabel metal1 12415 5202 12415 5202 0 net48
rlabel metal1 12323 3434 12323 3434 0 net49
rlabel metal2 1932 5236 1932 5236 0 net5
rlabel metal1 11239 5270 11239 5270 0 net50
rlabel metal1 3097 4182 3097 4182 0 net51
rlabel metal1 2724 4590 2724 4590 0 net52
rlabel metal1 3854 2414 3854 2414 0 net53
rlabel metal2 1610 9180 1610 9180 0 net6
rlabel metal1 1610 12240 1610 12240 0 net7
rlabel metal1 1610 13804 1610 13804 0 net8
rlabel metal1 1840 12206 1840 12206 0 net9
rlabel metal3 2384 2244 2384 2244 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 16000 20000
<< end >>
