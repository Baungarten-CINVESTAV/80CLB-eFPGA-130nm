// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype wire
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Feb  1 18:16:39 2024
//-------------------------------------------
// ----- Verilog module for fpga_top -----

//----- GLOBAL PORTS -----
wire prog_clk;
//----- GLOBAL PORTS -----
wire  set;
//----- GLOBAL PORTS -----
wire reset;
//----- GLOBAL PORTS -----
wire  clk;
//----- GPIO PORTS -----
wire [35:0] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
wire ccff_head;
//----- OUTPUT PORTS -----
wire ccff_tail;

assign prog_clk = io_in[36];
assign set = io_in[34];
assign reset = io_in[35];
assign clk = io_in[37];
assign {io_out[5],io_out[6],io_out[7],io_out[8],io_out[9],io_out[10],io_out[11]} = gfpga_pad_GPIO_PAD[19:13];
assign {io_out[14],io_out[15],io_out[16],io_out[17],io_out[18],io_out[19],io_out[20],io_out[21],io_out[22],io_out[23]} = gfpga_pad_GPIO_PAD[12:3];
assign gfpga_pad_GPIO_PAD[2:0] = {io_in[24],io_in[25],io_in[26]};
assign gfpga_pad_GPIO_PAD[35:29] = {io_in[27],io_in[28],io_in[29],io_in[30],io_in[31],io_in[32],io_in[33]};
assign ccff_head = io_in[12];
assign  io_out[13] = ccff_tail;
/*
assign io_oeb[21:19]={3{1'b1}}; // Inputs
assign io_oeb[28:22]={7{1'b1}}; // Inputs
assign  io_oeb[8:0]={9{1'b0}}; //Outputs
assign  io_oeb[18:9]={10{1'b0}}; //Outputs

assign io_oeb[37:29]={9{1'b0}}; // Inputs

assign  io_out[8:7]={2{1'b0}}; //Outputs
assign  io_out[37:19]=0; //Outputs
assign la_data_out = 128'b0;
*/

ioenb ioenb(
`ifdef USE_POWER_PINS
    .vccd1 (vccd1),	// User area 1 1.8V supply
    .vssd1 (vssd1),	// User area 1 digital ground
`endif
    .io_oeb (io_oeb)

);

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:8] cbx_1__0__0_chanx_left_out;
wire [0:8] cbx_1__0__0_chanx_right_out;
wire [0:8] cbx_1__0__1_chanx_left_out;
wire [0:8] cbx_1__0__1_chanx_right_out;
wire [0:8] cbx_1__0__2_chanx_left_out;
wire [0:8] cbx_1__0__2_chanx_right_out;
wire [0:8] cbx_1__0__3_chanx_left_out;
wire [0:8] cbx_1__0__3_chanx_right_out;
wire [0:8] cbx_1__0__4_chanx_left_out;
wire [0:8] cbx_1__0__4_chanx_right_out;
wire [0:8] cbx_1__0__5_chanx_left_out;
wire [0:8] cbx_1__0__5_chanx_right_out;
wire [0:8] cbx_1__0__6_chanx_left_out;
wire [0:8] cbx_1__0__6_chanx_right_out;
wire [0:8] cbx_1__0__7_chanx_left_out;
wire [0:8] cbx_1__0__7_chanx_right_out;
wire [0:8] cbx_1__10__0_chanx_left_out;
wire [0:8] cbx_1__10__0_chanx_right_out;
wire [0:8] cbx_1__10__1_chanx_left_out;
wire [0:8] cbx_1__10__1_chanx_right_out;
wire [0:8] cbx_1__10__2_chanx_left_out;
wire [0:8] cbx_1__10__2_chanx_right_out;
wire [0:8] cbx_1__10__3_chanx_left_out;
wire [0:8] cbx_1__10__3_chanx_right_out;
wire [0:8] cbx_1__10__4_chanx_left_out;
wire [0:8] cbx_1__10__4_chanx_right_out;
wire [0:8] cbx_1__10__5_chanx_left_out;
wire [0:8] cbx_1__10__5_chanx_right_out;
wire [0:8] cbx_1__10__6_chanx_left_out;
wire [0:8] cbx_1__10__6_chanx_right_out;
wire [0:8] cbx_1__10__7_chanx_left_out;
wire [0:8] cbx_1__10__7_chanx_right_out;
wire [0:8] cbx_1__1__0_chanx_left_out;
wire [0:8] cbx_1__1__0_chanx_right_out;
wire [0:8] cbx_1__1__10_chanx_left_out;
wire [0:8] cbx_1__1__10_chanx_right_out;
wire [0:8] cbx_1__1__11_chanx_left_out;
wire [0:8] cbx_1__1__11_chanx_right_out;
wire [0:8] cbx_1__1__12_chanx_left_out;
wire [0:8] cbx_1__1__12_chanx_right_out;
wire [0:8] cbx_1__1__13_chanx_left_out;
wire [0:8] cbx_1__1__13_chanx_right_out;
wire [0:8] cbx_1__1__14_chanx_left_out;
wire [0:8] cbx_1__1__14_chanx_right_out;
wire [0:8] cbx_1__1__15_chanx_left_out;
wire [0:8] cbx_1__1__15_chanx_right_out;
wire [0:8] cbx_1__1__16_chanx_left_out;
wire [0:8] cbx_1__1__16_chanx_right_out;
wire [0:8] cbx_1__1__17_chanx_left_out;
wire [0:8] cbx_1__1__17_chanx_right_out;
wire [0:8] cbx_1__1__18_chanx_left_out;
wire [0:8] cbx_1__1__18_chanx_right_out;
wire [0:8] cbx_1__1__19_chanx_left_out;
wire [0:8] cbx_1__1__19_chanx_right_out;
wire [0:8] cbx_1__1__1_chanx_left_out;
wire [0:8] cbx_1__1__1_chanx_right_out;
wire [0:8] cbx_1__1__20_chanx_left_out;
wire [0:8] cbx_1__1__20_chanx_right_out;
wire [0:8] cbx_1__1__21_chanx_left_out;
wire [0:8] cbx_1__1__21_chanx_right_out;
wire [0:8] cbx_1__1__22_chanx_left_out;
wire [0:8] cbx_1__1__22_chanx_right_out;
wire [0:8] cbx_1__1__23_chanx_left_out;
wire [0:8] cbx_1__1__23_chanx_right_out;
wire [0:8] cbx_1__1__24_chanx_left_out;
wire [0:8] cbx_1__1__24_chanx_right_out;
wire [0:8] cbx_1__1__25_chanx_left_out;
wire [0:8] cbx_1__1__25_chanx_right_out;
wire [0:8] cbx_1__1__26_chanx_left_out;
wire [0:8] cbx_1__1__26_chanx_right_out;
wire [0:8] cbx_1__1__27_chanx_left_out;
wire [0:8] cbx_1__1__27_chanx_right_out;
wire [0:8] cbx_1__1__28_chanx_left_out;
wire [0:8] cbx_1__1__28_chanx_right_out;
wire [0:8] cbx_1__1__29_chanx_left_out;
wire [0:8] cbx_1__1__29_chanx_right_out;
wire [0:8] cbx_1__1__2_chanx_left_out;
wire [0:8] cbx_1__1__2_chanx_right_out;
wire [0:8] cbx_1__1__30_chanx_left_out;
wire [0:8] cbx_1__1__30_chanx_right_out;
wire [0:8] cbx_1__1__31_chanx_left_out;
wire [0:8] cbx_1__1__31_chanx_right_out;
wire [0:8] cbx_1__1__32_chanx_left_out;
wire [0:8] cbx_1__1__32_chanx_right_out;
wire [0:8] cbx_1__1__33_chanx_left_out;
wire [0:8] cbx_1__1__33_chanx_right_out;
wire [0:8] cbx_1__1__34_chanx_left_out;
wire [0:8] cbx_1__1__34_chanx_right_out;
wire [0:8] cbx_1__1__35_chanx_left_out;
wire [0:8] cbx_1__1__35_chanx_right_out;
wire [0:8] cbx_1__1__36_chanx_left_out;
wire [0:8] cbx_1__1__36_chanx_right_out;
wire [0:8] cbx_1__1__37_chanx_left_out;
wire [0:8] cbx_1__1__37_chanx_right_out;
wire [0:8] cbx_1__1__38_chanx_left_out;
wire [0:8] cbx_1__1__38_chanx_right_out;
wire [0:8] cbx_1__1__39_chanx_left_out;
wire [0:8] cbx_1__1__39_chanx_right_out;
wire [0:8] cbx_1__1__3_chanx_left_out;
wire [0:8] cbx_1__1__3_chanx_right_out;
wire [0:8] cbx_1__1__40_chanx_left_out;
wire [0:8] cbx_1__1__40_chanx_right_out;
wire [0:8] cbx_1__1__41_chanx_left_out;
wire [0:8] cbx_1__1__41_chanx_right_out;
wire [0:8] cbx_1__1__42_chanx_left_out;
wire [0:8] cbx_1__1__42_chanx_right_out;
wire [0:8] cbx_1__1__43_chanx_left_out;
wire [0:8] cbx_1__1__43_chanx_right_out;
wire [0:8] cbx_1__1__44_chanx_left_out;
wire [0:8] cbx_1__1__44_chanx_right_out;
wire [0:8] cbx_1__1__45_chanx_left_out;
wire [0:8] cbx_1__1__45_chanx_right_out;
wire [0:8] cbx_1__1__46_chanx_left_out;
wire [0:8] cbx_1__1__46_chanx_right_out;
wire [0:8] cbx_1__1__47_chanx_left_out;
wire [0:8] cbx_1__1__47_chanx_right_out;
wire [0:8] cbx_1__1__48_chanx_left_out;
wire [0:8] cbx_1__1__48_chanx_right_out;
wire [0:8] cbx_1__1__49_chanx_left_out;
wire [0:8] cbx_1__1__49_chanx_right_out;
wire [0:8] cbx_1__1__4_chanx_left_out;
wire [0:8] cbx_1__1__4_chanx_right_out;
wire [0:8] cbx_1__1__50_chanx_left_out;
wire [0:8] cbx_1__1__50_chanx_right_out;
wire [0:8] cbx_1__1__51_chanx_left_out;
wire [0:8] cbx_1__1__51_chanx_right_out;
wire [0:8] cbx_1__1__52_chanx_left_out;
wire [0:8] cbx_1__1__52_chanx_right_out;
wire [0:8] cbx_1__1__53_chanx_left_out;
wire [0:8] cbx_1__1__53_chanx_right_out;
wire [0:8] cbx_1__1__54_chanx_left_out;
wire [0:8] cbx_1__1__54_chanx_right_out;
wire [0:8] cbx_1__1__55_chanx_left_out;
wire [0:8] cbx_1__1__55_chanx_right_out;
wire [0:8] cbx_1__1__56_chanx_left_out;
wire [0:8] cbx_1__1__56_chanx_right_out;
wire [0:8] cbx_1__1__57_chanx_left_out;
wire [0:8] cbx_1__1__57_chanx_right_out;
wire [0:8] cbx_1__1__58_chanx_left_out;
wire [0:8] cbx_1__1__58_chanx_right_out;
wire [0:8] cbx_1__1__59_chanx_left_out;
wire [0:8] cbx_1__1__59_chanx_right_out;
wire [0:8] cbx_1__1__5_chanx_left_out;
wire [0:8] cbx_1__1__5_chanx_right_out;
wire [0:8] cbx_1__1__60_chanx_left_out;
wire [0:8] cbx_1__1__60_chanx_right_out;
wire [0:8] cbx_1__1__61_chanx_left_out;
wire [0:8] cbx_1__1__61_chanx_right_out;
wire [0:8] cbx_1__1__62_chanx_left_out;
wire [0:8] cbx_1__1__62_chanx_right_out;
wire [0:8] cbx_1__1__63_chanx_left_out;
wire [0:8] cbx_1__1__63_chanx_right_out;
wire [0:8] cbx_1__1__64_chanx_left_out;
wire [0:8] cbx_1__1__64_chanx_right_out;
wire [0:8] cbx_1__1__65_chanx_left_out;
wire [0:8] cbx_1__1__65_chanx_right_out;
wire [0:8] cbx_1__1__66_chanx_left_out;
wire [0:8] cbx_1__1__66_chanx_right_out;
wire [0:8] cbx_1__1__67_chanx_left_out;
wire [0:8] cbx_1__1__67_chanx_right_out;
wire [0:8] cbx_1__1__68_chanx_left_out;
wire [0:8] cbx_1__1__68_chanx_right_out;
wire [0:8] cbx_1__1__69_chanx_left_out;
wire [0:8] cbx_1__1__69_chanx_right_out;
wire [0:8] cbx_1__1__6_chanx_left_out;
wire [0:8] cbx_1__1__6_chanx_right_out;
wire [0:8] cbx_1__1__70_chanx_left_out;
wire [0:8] cbx_1__1__70_chanx_right_out;
wire [0:8] cbx_1__1__71_chanx_left_out;
wire [0:8] cbx_1__1__71_chanx_right_out;
wire [0:8] cbx_1__1__7_chanx_left_out;
wire [0:8] cbx_1__1__7_chanx_right_out;
wire [0:8] cbx_1__1__8_chanx_left_out;
wire [0:8] cbx_1__1__8_chanx_right_out;
wire [0:8] cbx_1__1__9_chanx_left_out;
wire [0:8] cbx_1__1__9_chanx_right_out;
wire [0:8] cby_0__1__0_chany_bottom_out;
wire [0:8] cby_0__1__0_chany_top_out;
wire [0:8] cby_0__1__1_chany_bottom_out;
wire [0:8] cby_0__1__1_chany_top_out;
wire [0:8] cby_0__1__2_chany_bottom_out;
wire [0:8] cby_0__1__2_chany_top_out;
wire [0:8] cby_0__1__3_chany_bottom_out;
wire [0:8] cby_0__1__3_chany_top_out;
wire [0:8] cby_0__1__4_chany_bottom_out;
wire [0:8] cby_0__1__4_chany_top_out;
wire [0:8] cby_0__1__5_chany_bottom_out;
wire [0:8] cby_0__1__5_chany_top_out;
wire [0:8] cby_0__1__6_chany_bottom_out;
wire [0:8] cby_0__1__6_chany_top_out;
wire [0:8] cby_0__1__7_chany_bottom_out;
wire [0:8] cby_0__1__7_chany_top_out;
wire [0:8] cby_0__1__8_chany_bottom_out;
wire [0:8] cby_0__1__8_chany_top_out;
wire [0:8] cby_0__1__9_chany_bottom_out;
wire [0:8] cby_0__1__9_chany_top_out;
wire [0:8] cby_1__1__0_chany_bottom_out;
wire [0:8] cby_1__1__0_chany_top_out;
wire [0:8] cby_1__1__10_chany_bottom_out;
wire [0:8] cby_1__1__10_chany_top_out;
wire [0:8] cby_1__1__11_chany_bottom_out;
wire [0:8] cby_1__1__11_chany_top_out;
wire [0:8] cby_1__1__12_chany_bottom_out;
wire [0:8] cby_1__1__12_chany_top_out;
wire [0:8] cby_1__1__13_chany_bottom_out;
wire [0:8] cby_1__1__13_chany_top_out;
wire [0:8] cby_1__1__14_chany_bottom_out;
wire [0:8] cby_1__1__14_chany_top_out;
wire [0:8] cby_1__1__15_chany_bottom_out;
wire [0:8] cby_1__1__15_chany_top_out;
wire [0:8] cby_1__1__16_chany_bottom_out;
wire [0:8] cby_1__1__16_chany_top_out;
wire [0:8] cby_1__1__17_chany_bottom_out;
wire [0:8] cby_1__1__17_chany_top_out;
wire [0:8] cby_1__1__18_chany_bottom_out;
wire [0:8] cby_1__1__18_chany_top_out;
wire [0:8] cby_1__1__19_chany_bottom_out;
wire [0:8] cby_1__1__19_chany_top_out;
wire [0:8] cby_1__1__1_chany_bottom_out;
wire [0:8] cby_1__1__1_chany_top_out;
wire [0:8] cby_1__1__20_chany_bottom_out;
wire [0:8] cby_1__1__20_chany_top_out;
wire [0:8] cby_1__1__21_chany_bottom_out;
wire [0:8] cby_1__1__21_chany_top_out;
wire [0:8] cby_1__1__22_chany_bottom_out;
wire [0:8] cby_1__1__22_chany_top_out;
wire [0:8] cby_1__1__23_chany_bottom_out;
wire [0:8] cby_1__1__23_chany_top_out;
wire [0:8] cby_1__1__24_chany_bottom_out;
wire [0:8] cby_1__1__24_chany_top_out;
wire [0:8] cby_1__1__25_chany_bottom_out;
wire [0:8] cby_1__1__25_chany_top_out;
wire [0:8] cby_1__1__26_chany_bottom_out;
wire [0:8] cby_1__1__26_chany_top_out;
wire [0:8] cby_1__1__27_chany_bottom_out;
wire [0:8] cby_1__1__27_chany_top_out;
wire [0:8] cby_1__1__28_chany_bottom_out;
wire [0:8] cby_1__1__28_chany_top_out;
wire [0:8] cby_1__1__29_chany_bottom_out;
wire [0:8] cby_1__1__29_chany_top_out;
wire [0:8] cby_1__1__2_chany_bottom_out;
wire [0:8] cby_1__1__2_chany_top_out;
wire [0:8] cby_1__1__30_chany_bottom_out;
wire [0:8] cby_1__1__30_chany_top_out;
wire [0:8] cby_1__1__31_chany_bottom_out;
wire [0:8] cby_1__1__31_chany_top_out;
wire [0:8] cby_1__1__32_chany_bottom_out;
wire [0:8] cby_1__1__32_chany_top_out;
wire [0:8] cby_1__1__33_chany_bottom_out;
wire [0:8] cby_1__1__33_chany_top_out;
wire [0:8] cby_1__1__34_chany_bottom_out;
wire [0:8] cby_1__1__34_chany_top_out;
wire [0:8] cby_1__1__35_chany_bottom_out;
wire [0:8] cby_1__1__35_chany_top_out;
wire [0:8] cby_1__1__36_chany_bottom_out;
wire [0:8] cby_1__1__36_chany_top_out;
wire [0:8] cby_1__1__37_chany_bottom_out;
wire [0:8] cby_1__1__37_chany_top_out;
wire [0:8] cby_1__1__38_chany_bottom_out;
wire [0:8] cby_1__1__38_chany_top_out;
wire [0:8] cby_1__1__39_chany_bottom_out;
wire [0:8] cby_1__1__39_chany_top_out;
wire [0:8] cby_1__1__3_chany_bottom_out;
wire [0:8] cby_1__1__3_chany_top_out;
wire [0:8] cby_1__1__40_chany_bottom_out;
wire [0:8] cby_1__1__40_chany_top_out;
wire [0:8] cby_1__1__41_chany_bottom_out;
wire [0:8] cby_1__1__41_chany_top_out;
wire [0:8] cby_1__1__42_chany_bottom_out;
wire [0:8] cby_1__1__42_chany_top_out;
wire [0:8] cby_1__1__43_chany_bottom_out;
wire [0:8] cby_1__1__43_chany_top_out;
wire [0:8] cby_1__1__44_chany_bottom_out;
wire [0:8] cby_1__1__44_chany_top_out;
wire [0:8] cby_1__1__45_chany_bottom_out;
wire [0:8] cby_1__1__45_chany_top_out;
wire [0:8] cby_1__1__46_chany_bottom_out;
wire [0:8] cby_1__1__46_chany_top_out;
wire [0:8] cby_1__1__47_chany_bottom_out;
wire [0:8] cby_1__1__47_chany_top_out;
wire [0:8] cby_1__1__48_chany_bottom_out;
wire [0:8] cby_1__1__48_chany_top_out;
wire [0:8] cby_1__1__49_chany_bottom_out;
wire [0:8] cby_1__1__49_chany_top_out;
wire [0:8] cby_1__1__4_chany_bottom_out;
wire [0:8] cby_1__1__4_chany_top_out;
wire [0:8] cby_1__1__50_chany_bottom_out;
wire [0:8] cby_1__1__50_chany_top_out;
wire [0:8] cby_1__1__51_chany_bottom_out;
wire [0:8] cby_1__1__51_chany_top_out;
wire [0:8] cby_1__1__52_chany_bottom_out;
wire [0:8] cby_1__1__52_chany_top_out;
wire [0:8] cby_1__1__53_chany_bottom_out;
wire [0:8] cby_1__1__53_chany_top_out;
wire [0:8] cby_1__1__54_chany_bottom_out;
wire [0:8] cby_1__1__54_chany_top_out;
wire [0:8] cby_1__1__55_chany_bottom_out;
wire [0:8] cby_1__1__55_chany_top_out;
wire [0:8] cby_1__1__56_chany_bottom_out;
wire [0:8] cby_1__1__56_chany_top_out;
wire [0:8] cby_1__1__57_chany_bottom_out;
wire [0:8] cby_1__1__57_chany_top_out;
wire [0:8] cby_1__1__58_chany_bottom_out;
wire [0:8] cby_1__1__58_chany_top_out;
wire [0:8] cby_1__1__59_chany_bottom_out;
wire [0:8] cby_1__1__59_chany_top_out;
wire [0:8] cby_1__1__5_chany_bottom_out;
wire [0:8] cby_1__1__5_chany_top_out;
wire [0:8] cby_1__1__60_chany_bottom_out;
wire [0:8] cby_1__1__60_chany_top_out;
wire [0:8] cby_1__1__61_chany_bottom_out;
wire [0:8] cby_1__1__61_chany_top_out;
wire [0:8] cby_1__1__62_chany_bottom_out;
wire [0:8] cby_1__1__62_chany_top_out;
wire [0:8] cby_1__1__63_chany_bottom_out;
wire [0:8] cby_1__1__63_chany_top_out;
wire [0:8] cby_1__1__64_chany_bottom_out;
wire [0:8] cby_1__1__64_chany_top_out;
wire [0:8] cby_1__1__65_chany_bottom_out;
wire [0:8] cby_1__1__65_chany_top_out;
wire [0:8] cby_1__1__66_chany_bottom_out;
wire [0:8] cby_1__1__66_chany_top_out;
wire [0:8] cby_1__1__67_chany_bottom_out;
wire [0:8] cby_1__1__67_chany_top_out;
wire [0:8] cby_1__1__68_chany_bottom_out;
wire [0:8] cby_1__1__68_chany_top_out;
wire [0:8] cby_1__1__69_chany_bottom_out;
wire [0:8] cby_1__1__69_chany_top_out;
wire [0:8] cby_1__1__6_chany_bottom_out;
wire [0:8] cby_1__1__6_chany_top_out;
wire [0:8] cby_1__1__7_chany_bottom_out;
wire [0:8] cby_1__1__7_chany_top_out;
wire [0:8] cby_1__1__8_chany_bottom_out;
wire [0:8] cby_1__1__8_chany_top_out;
wire [0:8] cby_1__1__9_chany_bottom_out;
wire [0:8] cby_1__1__9_chany_top_out;
wire [0:8] cby_8__1__0_chany_bottom_out;
wire [0:8] cby_8__1__0_chany_top_out;
wire [0:8] cby_8__1__1_chany_bottom_out;
wire [0:8] cby_8__1__1_chany_top_out;
wire [0:8] cby_8__1__2_chany_bottom_out;
wire [0:8] cby_8__1__2_chany_top_out;
wire [0:8] cby_8__1__3_chany_bottom_out;
wire [0:8] cby_8__1__3_chany_top_out;
wire [0:8] cby_8__1__4_chany_bottom_out;
wire [0:8] cby_8__1__4_chany_top_out;
wire [0:8] cby_8__1__5_chany_bottom_out;
wire [0:8] cby_8__1__5_chany_top_out;
wire [0:8] cby_8__1__6_chany_bottom_out;
wire [0:8] cby_8__1__6_chany_top_out;
wire [0:8] cby_8__1__7_chany_bottom_out;
wire [0:8] cby_8__1__7_chany_top_out;
wire [0:8] cby_8__1__8_chany_bottom_out;
wire [0:8] cby_8__1__8_chany_top_out;
wire [0:8] cby_8__1__9_chany_bottom_out;
wire [0:8] cby_8__1__9_chany_top_out;
wire [0:8] sb_0__0__0_chanx_right_out;
wire [0:8] sb_0__0__0_chany_top_out;
wire [0:8] sb_0__10__0_chanx_right_out;
wire [0:8] sb_0__10__0_chany_bottom_out;
wire [0:8] sb_0__1__0_chanx_right_out;
wire [0:8] sb_0__1__0_chany_bottom_out;
wire [0:8] sb_0__1__0_chany_top_out;
wire [0:8] sb_0__1__1_chanx_right_out;
wire [0:8] sb_0__1__1_chany_bottom_out;
wire [0:8] sb_0__1__1_chany_top_out;
wire [0:8] sb_0__1__2_chanx_right_out;
wire [0:8] sb_0__1__2_chany_bottom_out;
wire [0:8] sb_0__1__2_chany_top_out;
wire [0:8] sb_0__1__3_chanx_right_out;
wire [0:8] sb_0__1__3_chany_bottom_out;
wire [0:8] sb_0__1__3_chany_top_out;
wire [0:8] sb_0__1__4_chanx_right_out;
wire [0:8] sb_0__1__4_chany_bottom_out;
wire [0:8] sb_0__1__4_chany_top_out;
wire [0:8] sb_0__1__5_chanx_right_out;
wire [0:8] sb_0__1__5_chany_bottom_out;
wire [0:8] sb_0__1__5_chany_top_out;
wire [0:8] sb_0__1__6_chanx_right_out;
wire [0:8] sb_0__1__6_chany_bottom_out;
wire [0:8] sb_0__1__6_chany_top_out;
wire [0:8] sb_0__1__7_chanx_right_out;
wire [0:8] sb_0__1__7_chany_bottom_out;
wire [0:8] sb_0__1__7_chany_top_out;
wire [0:8] sb_0__1__8_chanx_right_out;
wire [0:8] sb_0__1__8_chany_bottom_out;
wire [0:8] sb_0__1__8_chany_top_out;
wire [0:8] sb_1__0__0_chanx_left_out;
wire [0:8] sb_1__0__0_chanx_right_out;
wire [0:8] sb_1__0__0_chany_top_out;
wire [0:8] sb_1__0__1_chanx_left_out;
wire [0:8] sb_1__0__1_chanx_right_out;
wire [0:8] sb_1__0__1_chany_top_out;
wire [0:8] sb_1__0__2_chanx_left_out;
wire [0:8] sb_1__0__2_chanx_right_out;
wire [0:8] sb_1__0__2_chany_top_out;
wire [0:8] sb_1__0__3_chanx_left_out;
wire [0:8] sb_1__0__3_chanx_right_out;
wire [0:8] sb_1__0__3_chany_top_out;
wire [0:8] sb_1__0__4_chanx_left_out;
wire [0:8] sb_1__0__4_chanx_right_out;
wire [0:8] sb_1__0__4_chany_top_out;
wire [0:8] sb_1__0__5_chanx_left_out;
wire [0:8] sb_1__0__5_chanx_right_out;
wire [0:8] sb_1__0__5_chany_top_out;
wire [0:8] sb_1__0__6_chanx_left_out;
wire [0:8] sb_1__0__6_chanx_right_out;
wire [0:8] sb_1__0__6_chany_top_out;
wire [0:8] sb_1__10__0_chanx_left_out;
wire [0:8] sb_1__10__0_chanx_right_out;
wire [0:8] sb_1__10__0_chany_bottom_out;
wire [0:8] sb_1__10__1_chanx_left_out;
wire [0:8] sb_1__10__1_chanx_right_out;
wire [0:8] sb_1__10__1_chany_bottom_out;
wire [0:8] sb_1__10__2_chanx_left_out;
wire [0:8] sb_1__10__2_chanx_right_out;
wire [0:8] sb_1__10__2_chany_bottom_out;
wire [0:8] sb_1__10__3_chanx_left_out;
wire [0:8] sb_1__10__3_chanx_right_out;
wire [0:8] sb_1__10__3_chany_bottom_out;
wire [0:8] sb_1__10__4_chanx_left_out;
wire [0:8] sb_1__10__4_chanx_right_out;
wire [0:8] sb_1__10__4_chany_bottom_out;
wire [0:8] sb_1__10__5_chanx_left_out;
wire [0:8] sb_1__10__5_chanx_right_out;
wire [0:8] sb_1__10__5_chany_bottom_out;
wire [0:8] sb_1__10__6_chanx_left_out;
wire [0:8] sb_1__10__6_chanx_right_out;
wire [0:8] sb_1__10__6_chany_bottom_out;
wire [0:8] sb_1__1__0_chanx_left_out;
wire [0:8] sb_1__1__0_chanx_right_out;
wire [0:8] sb_1__1__0_chany_bottom_out;
wire [0:8] sb_1__1__0_chany_top_out;
wire [0:8] sb_1__1__10_chanx_left_out;
wire [0:8] sb_1__1__10_chanx_right_out;
wire [0:8] sb_1__1__10_chany_bottom_out;
wire [0:8] sb_1__1__10_chany_top_out;
wire [0:8] sb_1__1__11_chanx_left_out;
wire [0:8] sb_1__1__11_chanx_right_out;
wire [0:8] sb_1__1__11_chany_bottom_out;
wire [0:8] sb_1__1__11_chany_top_out;
wire [0:8] sb_1__1__12_chanx_left_out;
wire [0:8] sb_1__1__12_chanx_right_out;
wire [0:8] sb_1__1__12_chany_bottom_out;
wire [0:8] sb_1__1__12_chany_top_out;
wire [0:8] sb_1__1__13_chanx_left_out;
wire [0:8] sb_1__1__13_chanx_right_out;
wire [0:8] sb_1__1__13_chany_bottom_out;
wire [0:8] sb_1__1__13_chany_top_out;
wire [0:8] sb_1__1__14_chanx_left_out;
wire [0:8] sb_1__1__14_chanx_right_out;
wire [0:8] sb_1__1__14_chany_bottom_out;
wire [0:8] sb_1__1__14_chany_top_out;
wire [0:8] sb_1__1__15_chanx_left_out;
wire [0:8] sb_1__1__15_chanx_right_out;
wire [0:8] sb_1__1__15_chany_bottom_out;
wire [0:8] sb_1__1__15_chany_top_out;
wire [0:8] sb_1__1__16_chanx_left_out;
wire [0:8] sb_1__1__16_chanx_right_out;
wire [0:8] sb_1__1__16_chany_bottom_out;
wire [0:8] sb_1__1__16_chany_top_out;
wire [0:8] sb_1__1__17_chanx_left_out;
wire [0:8] sb_1__1__17_chanx_right_out;
wire [0:8] sb_1__1__17_chany_bottom_out;
wire [0:8] sb_1__1__17_chany_top_out;
wire [0:8] sb_1__1__18_chanx_left_out;
wire [0:8] sb_1__1__18_chanx_right_out;
wire [0:8] sb_1__1__18_chany_bottom_out;
wire [0:8] sb_1__1__18_chany_top_out;
wire [0:8] sb_1__1__19_chanx_left_out;
wire [0:8] sb_1__1__19_chanx_right_out;
wire [0:8] sb_1__1__19_chany_bottom_out;
wire [0:8] sb_1__1__19_chany_top_out;
wire [0:8] sb_1__1__1_chanx_left_out;
wire [0:8] sb_1__1__1_chanx_right_out;
wire [0:8] sb_1__1__1_chany_bottom_out;
wire [0:8] sb_1__1__1_chany_top_out;
wire [0:8] sb_1__1__20_chanx_left_out;
wire [0:8] sb_1__1__20_chanx_right_out;
wire [0:8] sb_1__1__20_chany_bottom_out;
wire [0:8] sb_1__1__20_chany_top_out;
wire [0:8] sb_1__1__21_chanx_left_out;
wire [0:8] sb_1__1__21_chanx_right_out;
wire [0:8] sb_1__1__21_chany_bottom_out;
wire [0:8] sb_1__1__21_chany_top_out;
wire [0:8] sb_1__1__22_chanx_left_out;
wire [0:8] sb_1__1__22_chanx_right_out;
wire [0:8] sb_1__1__22_chany_bottom_out;
wire [0:8] sb_1__1__22_chany_top_out;
wire [0:8] sb_1__1__23_chanx_left_out;
wire [0:8] sb_1__1__23_chanx_right_out;
wire [0:8] sb_1__1__23_chany_bottom_out;
wire [0:8] sb_1__1__23_chany_top_out;
wire [0:8] sb_1__1__24_chanx_left_out;
wire [0:8] sb_1__1__24_chanx_right_out;
wire [0:8] sb_1__1__24_chany_bottom_out;
wire [0:8] sb_1__1__24_chany_top_out;
wire [0:8] sb_1__1__25_chanx_left_out;
wire [0:8] sb_1__1__25_chanx_right_out;
wire [0:8] sb_1__1__25_chany_bottom_out;
wire [0:8] sb_1__1__25_chany_top_out;
wire [0:8] sb_1__1__26_chanx_left_out;
wire [0:8] sb_1__1__26_chanx_right_out;
wire [0:8] sb_1__1__26_chany_bottom_out;
wire [0:8] sb_1__1__26_chany_top_out;
wire [0:8] sb_1__1__27_chanx_left_out;
wire [0:8] sb_1__1__27_chanx_right_out;
wire [0:8] sb_1__1__27_chany_bottom_out;
wire [0:8] sb_1__1__27_chany_top_out;
wire [0:8] sb_1__1__28_chanx_left_out;
wire [0:8] sb_1__1__28_chanx_right_out;
wire [0:8] sb_1__1__28_chany_bottom_out;
wire [0:8] sb_1__1__28_chany_top_out;
wire [0:8] sb_1__1__29_chanx_left_out;
wire [0:8] sb_1__1__29_chanx_right_out;
wire [0:8] sb_1__1__29_chany_bottom_out;
wire [0:8] sb_1__1__29_chany_top_out;
wire [0:8] sb_1__1__2_chanx_left_out;
wire [0:8] sb_1__1__2_chanx_right_out;
wire [0:8] sb_1__1__2_chany_bottom_out;
wire [0:8] sb_1__1__2_chany_top_out;
wire [0:8] sb_1__1__30_chanx_left_out;
wire [0:8] sb_1__1__30_chanx_right_out;
wire [0:8] sb_1__1__30_chany_bottom_out;
wire [0:8] sb_1__1__30_chany_top_out;
wire [0:8] sb_1__1__31_chanx_left_out;
wire [0:8] sb_1__1__31_chanx_right_out;
wire [0:8] sb_1__1__31_chany_bottom_out;
wire [0:8] sb_1__1__31_chany_top_out;
wire [0:8] sb_1__1__32_chanx_left_out;
wire [0:8] sb_1__1__32_chanx_right_out;
wire [0:8] sb_1__1__32_chany_bottom_out;
wire [0:8] sb_1__1__32_chany_top_out;
wire [0:8] sb_1__1__33_chanx_left_out;
wire [0:8] sb_1__1__33_chanx_right_out;
wire [0:8] sb_1__1__33_chany_bottom_out;
wire [0:8] sb_1__1__33_chany_top_out;
wire [0:8] sb_1__1__34_chanx_left_out;
wire [0:8] sb_1__1__34_chanx_right_out;
wire [0:8] sb_1__1__34_chany_bottom_out;
wire [0:8] sb_1__1__34_chany_top_out;
wire [0:8] sb_1__1__35_chanx_left_out;
wire [0:8] sb_1__1__35_chanx_right_out;
wire [0:8] sb_1__1__35_chany_bottom_out;
wire [0:8] sb_1__1__35_chany_top_out;
wire [0:8] sb_1__1__36_chanx_left_out;
wire [0:8] sb_1__1__36_chanx_right_out;
wire [0:8] sb_1__1__36_chany_bottom_out;
wire [0:8] sb_1__1__36_chany_top_out;
wire [0:8] sb_1__1__37_chanx_left_out;
wire [0:8] sb_1__1__37_chanx_right_out;
wire [0:8] sb_1__1__37_chany_bottom_out;
wire [0:8] sb_1__1__37_chany_top_out;
wire [0:8] sb_1__1__38_chanx_left_out;
wire [0:8] sb_1__1__38_chanx_right_out;
wire [0:8] sb_1__1__38_chany_bottom_out;
wire [0:8] sb_1__1__38_chany_top_out;
wire [0:8] sb_1__1__39_chanx_left_out;
wire [0:8] sb_1__1__39_chanx_right_out;
wire [0:8] sb_1__1__39_chany_bottom_out;
wire [0:8] sb_1__1__39_chany_top_out;
wire [0:8] sb_1__1__3_chanx_left_out;
wire [0:8] sb_1__1__3_chanx_right_out;
wire [0:8] sb_1__1__3_chany_bottom_out;
wire [0:8] sb_1__1__3_chany_top_out;
wire [0:8] sb_1__1__40_chanx_left_out;
wire [0:8] sb_1__1__40_chanx_right_out;
wire [0:8] sb_1__1__40_chany_bottom_out;
wire [0:8] sb_1__1__40_chany_top_out;
wire [0:8] sb_1__1__41_chanx_left_out;
wire [0:8] sb_1__1__41_chanx_right_out;
wire [0:8] sb_1__1__41_chany_bottom_out;
wire [0:8] sb_1__1__41_chany_top_out;
wire [0:8] sb_1__1__42_chanx_left_out;
wire [0:8] sb_1__1__42_chanx_right_out;
wire [0:8] sb_1__1__42_chany_bottom_out;
wire [0:8] sb_1__1__42_chany_top_out;
wire [0:8] sb_1__1__43_chanx_left_out;
wire [0:8] sb_1__1__43_chanx_right_out;
wire [0:8] sb_1__1__43_chany_bottom_out;
wire [0:8] sb_1__1__43_chany_top_out;
wire [0:8] sb_1__1__44_chanx_left_out;
wire [0:8] sb_1__1__44_chanx_right_out;
wire [0:8] sb_1__1__44_chany_bottom_out;
wire [0:8] sb_1__1__44_chany_top_out;
wire [0:8] sb_1__1__45_chanx_left_out;
wire [0:8] sb_1__1__45_chanx_right_out;
wire [0:8] sb_1__1__45_chany_bottom_out;
wire [0:8] sb_1__1__45_chany_top_out;
wire [0:8] sb_1__1__46_chanx_left_out;
wire [0:8] sb_1__1__46_chanx_right_out;
wire [0:8] sb_1__1__46_chany_bottom_out;
wire [0:8] sb_1__1__46_chany_top_out;
wire [0:8] sb_1__1__47_chanx_left_out;
wire [0:8] sb_1__1__47_chanx_right_out;
wire [0:8] sb_1__1__47_chany_bottom_out;
wire [0:8] sb_1__1__47_chany_top_out;
wire [0:8] sb_1__1__48_chanx_left_out;
wire [0:8] sb_1__1__48_chanx_right_out;
wire [0:8] sb_1__1__48_chany_bottom_out;
wire [0:8] sb_1__1__48_chany_top_out;
wire [0:8] sb_1__1__49_chanx_left_out;
wire [0:8] sb_1__1__49_chanx_right_out;
wire [0:8] sb_1__1__49_chany_bottom_out;
wire [0:8] sb_1__1__49_chany_top_out;
wire [0:8] sb_1__1__4_chanx_left_out;
wire [0:8] sb_1__1__4_chanx_right_out;
wire [0:8] sb_1__1__4_chany_bottom_out;
wire [0:8] sb_1__1__4_chany_top_out;
wire [0:8] sb_1__1__50_chanx_left_out;
wire [0:8] sb_1__1__50_chanx_right_out;
wire [0:8] sb_1__1__50_chany_bottom_out;
wire [0:8] sb_1__1__50_chany_top_out;
wire [0:8] sb_1__1__51_chanx_left_out;
wire [0:8] sb_1__1__51_chanx_right_out;
wire [0:8] sb_1__1__51_chany_bottom_out;
wire [0:8] sb_1__1__51_chany_top_out;
wire [0:8] sb_1__1__52_chanx_left_out;
wire [0:8] sb_1__1__52_chanx_right_out;
wire [0:8] sb_1__1__52_chany_bottom_out;
wire [0:8] sb_1__1__52_chany_top_out;
wire [0:8] sb_1__1__53_chanx_left_out;
wire [0:8] sb_1__1__53_chanx_right_out;
wire [0:8] sb_1__1__53_chany_bottom_out;
wire [0:8] sb_1__1__53_chany_top_out;
wire [0:8] sb_1__1__54_chanx_left_out;
wire [0:8] sb_1__1__54_chanx_right_out;
wire [0:8] sb_1__1__54_chany_bottom_out;
wire [0:8] sb_1__1__54_chany_top_out;
wire [0:8] sb_1__1__55_chanx_left_out;
wire [0:8] sb_1__1__55_chanx_right_out;
wire [0:8] sb_1__1__55_chany_bottom_out;
wire [0:8] sb_1__1__55_chany_top_out;
wire [0:8] sb_1__1__56_chanx_left_out;
wire [0:8] sb_1__1__56_chanx_right_out;
wire [0:8] sb_1__1__56_chany_bottom_out;
wire [0:8] sb_1__1__56_chany_top_out;
wire [0:8] sb_1__1__57_chanx_left_out;
wire [0:8] sb_1__1__57_chanx_right_out;
wire [0:8] sb_1__1__57_chany_bottom_out;
wire [0:8] sb_1__1__57_chany_top_out;
wire [0:8] sb_1__1__58_chanx_left_out;
wire [0:8] sb_1__1__58_chanx_right_out;
wire [0:8] sb_1__1__58_chany_bottom_out;
wire [0:8] sb_1__1__58_chany_top_out;
wire [0:8] sb_1__1__59_chanx_left_out;
wire [0:8] sb_1__1__59_chanx_right_out;
wire [0:8] sb_1__1__59_chany_bottom_out;
wire [0:8] sb_1__1__59_chany_top_out;
wire [0:8] sb_1__1__5_chanx_left_out;
wire [0:8] sb_1__1__5_chanx_right_out;
wire [0:8] sb_1__1__5_chany_bottom_out;
wire [0:8] sb_1__1__5_chany_top_out;
wire [0:8] sb_1__1__60_chanx_left_out;
wire [0:8] sb_1__1__60_chanx_right_out;
wire [0:8] sb_1__1__60_chany_bottom_out;
wire [0:8] sb_1__1__60_chany_top_out;
wire [0:8] sb_1__1__61_chanx_left_out;
wire [0:8] sb_1__1__61_chanx_right_out;
wire [0:8] sb_1__1__61_chany_bottom_out;
wire [0:8] sb_1__1__61_chany_top_out;
wire [0:8] sb_1__1__62_chanx_left_out;
wire [0:8] sb_1__1__62_chanx_right_out;
wire [0:8] sb_1__1__62_chany_bottom_out;
wire [0:8] sb_1__1__62_chany_top_out;
wire [0:8] sb_1__1__6_chanx_left_out;
wire [0:8] sb_1__1__6_chanx_right_out;
wire [0:8] sb_1__1__6_chany_bottom_out;
wire [0:8] sb_1__1__6_chany_top_out;
wire [0:8] sb_1__1__7_chanx_left_out;
wire [0:8] sb_1__1__7_chanx_right_out;
wire [0:8] sb_1__1__7_chany_bottom_out;
wire [0:8] sb_1__1__7_chany_top_out;
wire [0:8] sb_1__1__8_chanx_left_out;
wire [0:8] sb_1__1__8_chanx_right_out;
wire [0:8] sb_1__1__8_chany_bottom_out;
wire [0:8] sb_1__1__8_chany_top_out;
wire [0:8] sb_1__1__9_chanx_left_out;
wire [0:8] sb_1__1__9_chanx_right_out;
wire [0:8] sb_1__1__9_chany_bottom_out;
wire [0:8] sb_1__1__9_chany_top_out;
wire [0:8] sb_8__0__0_chanx_left_out;
wire [0:8] sb_8__0__0_chany_top_out;
wire [0:8] sb_8__10__0_chanx_left_out;
wire [0:8] sb_8__10__0_chany_bottom_out;
wire [0:8] sb_8__1__0_chanx_left_out;
wire [0:8] sb_8__1__0_chany_bottom_out;
wire [0:8] sb_8__1__0_chany_top_out;
wire [0:8] sb_8__1__1_chanx_left_out;
wire [0:8] sb_8__1__1_chany_bottom_out;
wire [0:8] sb_8__1__1_chany_top_out;
wire [0:8] sb_8__1__2_chanx_left_out;
wire [0:8] sb_8__1__2_chany_bottom_out;
wire [0:8] sb_8__1__2_chany_top_out;
wire [0:8] sb_8__1__3_chanx_left_out;
wire [0:8] sb_8__1__3_chany_bottom_out;
wire [0:8] sb_8__1__3_chany_top_out;
wire [0:8] sb_8__1__4_chanx_left_out;
wire [0:8] sb_8__1__4_chany_bottom_out;
wire [0:8] sb_8__1__4_chany_top_out;
wire [0:8] sb_8__1__5_chanx_left_out;
wire [0:8] sb_8__1__5_chany_bottom_out;
wire [0:8] sb_8__1__5_chany_top_out;
wire [0:8] sb_8__1__6_chanx_left_out;
wire [0:8] sb_8__1__6_chany_bottom_out;
wire [0:8] sb_8__1__6_chany_top_out;
wire [0:8] sb_8__1__7_chanx_left_out;
wire [0:8] sb_8__1__7_chany_bottom_out;
wire [0:8] sb_8__1__7_chany_top_out;
wire [0:8] sb_8__1__8_chanx_left_out;
wire [0:8] sb_8__1__8_chany_bottom_out;
wire [0:8] sb_8__1__8_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[1]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[2]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top_out grid_io_top_4__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[3]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_top_out grid_io_top_5__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[4]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_4_ccff_tail));

	grid_io_top_out grid_io_top_6__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[5]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_5_ccff_tail));

	grid_io_top_out grid_io_top_7__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[6]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__6_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_6_ccff_tail));

	grid_io_top_out grid_io_top_8__11_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cbx_1__10__7_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_top_7_ccff_tail));

	grid_io_right_out grid_io_right_9__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right_out grid_io_right_9__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[9]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right_out grid_io_right_9__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[10]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right_out grid_io_right_9__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[11]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right_out grid_io_right_9__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[12]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right_out grid_io_right_9__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[13]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_right_out grid_io_right_9__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[14]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_6_ccff_tail));

	grid_io_right_out grid_io_right_9__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[15]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_8_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_7_ccff_tail));

	grid_io_right_out grid_io_right_9__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_right_9_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_8_ccff_tail));

	grid_io_right_out grid_io_right_9__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[17]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_right_9_ccff_tail));

	grid_io_bottom_out grid_io_bottom_8__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[18]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom_out grid_io_bottom_7__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[19]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_6__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[20]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_5__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[21]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[22]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_4_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[23]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_5_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(grid_io_bottom_7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_6_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[25]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_7_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[26]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[27]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[28]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[29]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[30]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[31]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_io_left grid_io_left_0__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_6_ccff_tail));

	grid_io_left grid_io_left_0__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[33]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_7_ccff_tail));

	grid_io_left grid_io_left_0__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[34]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__8_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_8_ccff_tail));

	grid_io_left grid_io_left_0__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[35]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(cby_0__1__9_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_tail(grid_io_left_9_ccff_tail));

	grid_clb grid_clb_1__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_1__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_1__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_1__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_1__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_1__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_1__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_2__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_2__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_2__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_2__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_2__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_2__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_2__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_2__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_2__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_3__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_3__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_3__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__22_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_3__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__23_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_3__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__24_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_24_ccff_tail));

	grid_clb grid_clb_3__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__25_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_25_ccff_tail));

	grid_clb grid_clb_3__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__26_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_26_ccff_tail));

	grid_clb grid_clb_3__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__27_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_27_ccff_tail));

	grid_clb grid_clb_3__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__28_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_28_ccff_tail));

	grid_clb grid_clb_3__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__29_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_29_ccff_tail));

	grid_clb grid_clb_4__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__30_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_30_ccff_tail));

	grid_clb grid_clb_4__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__21_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__21_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__31_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_31_ccff_tail));

	grid_clb grid_clb_4__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__22_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__22_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__32_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_32_ccff_tail));

	grid_clb grid_clb_4__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__23_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__23_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__33_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_33_ccff_tail));

	grid_clb grid_clb_4__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__24_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__24_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__34_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_34_ccff_tail));

	grid_clb grid_clb_4__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__25_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__25_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__35_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_35_ccff_tail));

	grid_clb grid_clb_4__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__26_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__26_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__36_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_36_ccff_tail));

	grid_clb grid_clb_4__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__27_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__27_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__37_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_37_ccff_tail));

	grid_clb grid_clb_4__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__28_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__28_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__38_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_38_ccff_tail));

	grid_clb grid_clb_4__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__29_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__29_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__39_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_39_ccff_tail));

	grid_clb grid_clb_5__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__30_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__30_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__40_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_40_ccff_tail));

	grid_clb grid_clb_5__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__31_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__31_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__41_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_41_ccff_tail));

	grid_clb grid_clb_5__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__32_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__32_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__42_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_42_ccff_tail));

	grid_clb grid_clb_5__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__33_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__33_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__43_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_43_ccff_tail));

	grid_clb grid_clb_5__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__34_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__34_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__44_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_44_ccff_tail));

	grid_clb grid_clb_5__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__35_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__35_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__45_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_45_ccff_tail));

	grid_clb grid_clb_5__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__36_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__36_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__46_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_46_ccff_tail));

	grid_clb grid_clb_5__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__37_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__37_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__47_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_47_ccff_tail));

	grid_clb grid_clb_5__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__38_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__38_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__48_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_48_ccff_tail));

	grid_clb grid_clb_5__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__39_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__39_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__49_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_49_ccff_tail));

	grid_clb grid_clb_6__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__40_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__40_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__50_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_50_ccff_tail));

	grid_clb grid_clb_6__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__41_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__41_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__51_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_51_ccff_tail));

	grid_clb grid_clb_6__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__42_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__42_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__52_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_52_ccff_tail));

	grid_clb grid_clb_6__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__43_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__43_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__53_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_53_ccff_tail));

	grid_clb grid_clb_6__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__44_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__44_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__54_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_54_ccff_tail));

	grid_clb grid_clb_6__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__45_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__45_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__55_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_55_ccff_tail));

	grid_clb grid_clb_6__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__46_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__46_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__56_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_56_ccff_tail));

	grid_clb grid_clb_6__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__47_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__47_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__57_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_57_ccff_tail));

	grid_clb grid_clb_6__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__48_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__48_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__58_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_58_ccff_tail));

	grid_clb grid_clb_6__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__49_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__49_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__59_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_59_ccff_tail));

	grid_clb grid_clb_7__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__50_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__50_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__60_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_60_ccff_tail));

	grid_clb grid_clb_7__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__51_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__51_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__61_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_61_ccff_tail));

	grid_clb grid_clb_7__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__52_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__52_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__62_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_62_ccff_tail));

	grid_clb grid_clb_7__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__53_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__53_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__63_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_63_ccff_tail));

	grid_clb grid_clb_7__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__54_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__54_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__64_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_64_ccff_tail));

	grid_clb grid_clb_7__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__55_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__55_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__65_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_65_ccff_tail));

	grid_clb grid_clb_7__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__56_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__56_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__66_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_66_ccff_tail));

	grid_clb grid_clb_7__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__57_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__57_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__67_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_67_ccff_tail));

	grid_clb grid_clb_7__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__58_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__58_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__68_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_68_ccff_tail));

	grid_clb grid_clb_7__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__59_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__59_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__69_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_69_ccff_tail));

	grid_clb grid_clb_8__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__60_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__60_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_70_ccff_tail));

	grid_clb grid_clb_8__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__61_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__61_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_71_ccff_tail));

	grid_clb grid_clb_8__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__62_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__62_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_72_ccff_tail));

	grid_clb grid_clb_8__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__63_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__63_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_73_ccff_tail));

	grid_clb grid_clb_8__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__64_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__64_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_74_ccff_tail));

	grid_clb grid_clb_8__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__65_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__65_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_75_ccff_tail));

	grid_clb grid_clb_8__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__66_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__66_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_76_ccff_tail));

	grid_clb grid_clb_8__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__67_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__67_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_77_ccff_tail));

	grid_clb grid_clb_8__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__68_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__68_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_78_ccff_tail));

	grid_clb grid_clb_8__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__69_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__69_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_8__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_79_ccff_tail));

	sb_0__0_ sb_0__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:8]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:8]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__3_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__4_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__1_ sb_0__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__5_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_6_ccff_tail),
		.chany_top_out(sb_0__1__4_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__4_ccff_tail));

	sb_0__1_ sb_0__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__6_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_7_ccff_tail),
		.chany_top_out(sb_0__1__5_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__5_ccff_tail));

	sb_0__1_ sb_0__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__7_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_8_ccff_tail),
		.chany_top_out(sb_0__1__6_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__6_ccff_tail));

	sb_0__1_ sb_0__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__8_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_9_ccff_tail),
		.chany_top_out(sb_0__1__7_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__7_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__7_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__7_ccff_tail));

	sb_0__1_ sb_0__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_0__1__9_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(sb_0__10__0_ccff_tail),
		.chany_top_out(sb_0__1__8_chany_top_out[0:8]),
		.chanx_right_out(sb_0__1__8_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__1__8_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__1__8_ccff_tail));

	sb_0__10_ sb_0__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__0_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__10__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_0__10__0_chany_bottom_out[0:8]),
		.ccff_tail(sb_0__10__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__10_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__20_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__30_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_5__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__40_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_30_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__0_ sb_6__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__50_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_40_ccff_tail),
		.chany_top_out(sb_1__0__5_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__5_ccff_tail));

	sb_1__0_ sb_7__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__60_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_50_ccff_tail),
		.chany_top_out(sb_1__0__6_chany_top_out[0:8]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:8]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:8]),
		.ccff_tail(sb_1__0__6_ccff_tail));

	sb_1__1_ sb_1__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__3_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_1__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__4_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_1__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__5_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_1__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__6_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_1__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__7_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_1__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__8_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_1__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__9_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__1_ sb_2__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__11_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_1__1__9_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__9_ccff_tail));

	sb_1__1_ sb_2__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__12_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__10_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__10_ccff_tail));

	sb_1__1_ sb_2__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__13_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__20_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_1__1__11_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__11_ccff_tail));

	sb_1__1_ sb_2__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__14_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__21_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__1__12_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__12_ccff_tail));

	sb_1__1_ sb_2__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__15_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__22_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_25_ccff_tail),
		.chany_top_out(sb_1__1__13_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__13_ccff_tail));

	sb_1__1_ sb_2__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__16_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__23_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__1__14_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__14_ccff_tail));

	sb_1__1_ sb_2__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__17_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__24_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_27_ccff_tail),
		.chany_top_out(sb_1__1__15_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__15_ccff_tail));

	sb_1__1_ sb_2__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__18_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__25_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__1__16_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__16_ccff_tail));

	sb_1__1_ sb_2__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__19_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__26_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_29_ccff_tail),
		.chany_top_out(sb_1__1__17_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__17_ccff_tail));

	sb_1__1_ sb_3__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__21_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__27_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_31_ccff_tail),
		.chany_top_out(sb_1__1__18_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__18_ccff_tail));

	sb_1__1_ sb_3__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__22_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__28_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__1__19_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__19_ccff_tail));

	sb_1__1_ sb_3__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__23_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__29_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__20_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_33_ccff_tail),
		.chany_top_out(sb_1__1__20_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__20_ccff_tail));

	sb_1__1_ sb_3__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__24_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__30_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__21_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__1__21_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__21_ccff_tail));

	sb_1__1_ sb_3__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__25_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__31_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__22_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_35_ccff_tail),
		.chany_top_out(sb_1__1__22_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__22_ccff_tail));

	sb_1__1_ sb_3__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__26_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__32_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__23_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__1__23_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__23_ccff_tail));

	sb_1__1_ sb_3__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__27_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__33_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__24_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_37_ccff_tail),
		.chany_top_out(sb_1__1__24_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__24_ccff_tail));

	sb_1__1_ sb_3__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__28_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__34_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__25_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__1__25_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__25_ccff_tail));

	sb_1__1_ sb_3__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__29_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__35_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__26_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_39_ccff_tail),
		.chany_top_out(sb_1__1__26_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__26_ccff_tail));

	sb_1__1_ sb_4__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__31_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__36_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__27_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_41_ccff_tail),
		.chany_top_out(sb_1__1__27_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__27_ccff_tail));

	sb_1__1_ sb_4__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__32_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__37_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__28_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_1__1__28_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__28_ccff_tail));

	sb_1__1_ sb_4__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__33_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__38_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__29_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_43_ccff_tail),
		.chany_top_out(sb_1__1__29_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__29_ccff_tail));

	sb_1__1_ sb_4__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__34_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__39_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__30_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_24_ccff_tail),
		.chany_top_out(sb_1__1__30_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__30_ccff_tail));

	sb_1__1_ sb_4__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__35_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__40_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__31_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_45_ccff_tail),
		.chany_top_out(sb_1__1__31_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__31_ccff_tail));

	sb_1__1_ sb_4__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__36_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__41_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__32_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_26_ccff_tail),
		.chany_top_out(sb_1__1__32_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__32_ccff_tail));

	sb_1__1_ sb_4__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__37_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__42_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__33_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_47_ccff_tail),
		.chany_top_out(sb_1__1__33_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__33_ccff_tail));

	sb_1__1_ sb_4__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__38_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__43_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__34_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_28_ccff_tail),
		.chany_top_out(sb_1__1__34_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__34_ccff_tail));

	sb_1__1_ sb_4__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__39_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__44_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__35_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_49_ccff_tail),
		.chany_top_out(sb_1__1__35_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__35_ccff_tail));

	sb_1__1_ sb_5__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__41_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__45_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__36_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_51_ccff_tail),
		.chany_top_out(sb_1__1__36_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__36_ccff_tail));

	sb_1__1_ sb_5__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__42_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__46_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__37_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_32_ccff_tail),
		.chany_top_out(sb_1__1__37_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__37_ccff_tail));

	sb_1__1_ sb_5__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__43_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__47_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__38_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_53_ccff_tail),
		.chany_top_out(sb_1__1__38_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__38_ccff_tail));

	sb_1__1_ sb_5__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__44_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__48_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__39_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_34_ccff_tail),
		.chany_top_out(sb_1__1__39_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__39_ccff_tail));

	sb_1__1_ sb_5__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__45_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__49_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__40_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_55_ccff_tail),
		.chany_top_out(sb_1__1__40_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__40_ccff_tail));

	sb_1__1_ sb_5__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__46_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__50_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__41_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_36_ccff_tail),
		.chany_top_out(sb_1__1__41_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__41_ccff_tail));

	sb_1__1_ sb_5__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__47_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__51_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__42_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_57_ccff_tail),
		.chany_top_out(sb_1__1__42_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__42_ccff_tail));

	sb_1__1_ sb_5__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__48_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__52_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__43_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_38_ccff_tail),
		.chany_top_out(sb_1__1__43_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__43_ccff_tail));

	sb_1__1_ sb_5__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__49_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__53_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__44_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_59_ccff_tail),
		.chany_top_out(sb_1__1__44_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__44_ccff_tail));

	sb_1__1_ sb_6__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__51_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__54_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__45_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_61_ccff_tail),
		.chany_top_out(sb_1__1__45_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__45_ccff_tail));

	sb_1__1_ sb_6__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__52_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__55_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__46_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_42_ccff_tail),
		.chany_top_out(sb_1__1__46_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__46_ccff_tail));

	sb_1__1_ sb_6__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__53_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__56_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__47_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_63_ccff_tail),
		.chany_top_out(sb_1__1__47_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__47_ccff_tail));

	sb_1__1_ sb_6__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__54_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__57_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__48_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_44_ccff_tail),
		.chany_top_out(sb_1__1__48_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__48_ccff_tail));

	sb_1__1_ sb_6__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__55_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__58_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__49_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_65_ccff_tail),
		.chany_top_out(sb_1__1__49_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__49_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__49_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__49_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__49_ccff_tail));

	sb_1__1_ sb_6__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__56_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__59_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__50_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_46_ccff_tail),
		.chany_top_out(sb_1__1__50_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__50_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__50_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__50_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__50_ccff_tail));

	sb_1__1_ sb_6__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__57_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__60_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__56_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__51_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_67_ccff_tail),
		.chany_top_out(sb_1__1__51_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__51_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__51_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__51_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__51_ccff_tail));

	sb_1__1_ sb_6__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__58_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__61_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__57_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__52_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_48_ccff_tail),
		.chany_top_out(sb_1__1__52_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__52_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__52_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__52_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__52_ccff_tail));

	sb_1__1_ sb_6__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__59_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__62_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__58_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__53_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_69_ccff_tail),
		.chany_top_out(sb_1__1__53_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__53_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__53_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__53_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__53_ccff_tail));

	sb_1__1_ sb_7__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__61_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__63_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__60_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__54_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_71_ccff_tail),
		.chany_top_out(sb_1__1__54_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__54_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__54_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__54_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__54_ccff_tail));

	sb_1__1_ sb_7__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__62_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__64_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__61_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__55_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_52_ccff_tail),
		.chany_top_out(sb_1__1__55_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__55_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__55_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__55_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__55_ccff_tail));

	sb_1__1_ sb_7__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__63_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__65_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__62_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__56_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_73_ccff_tail),
		.chany_top_out(sb_1__1__56_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__56_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__56_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__56_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__56_ccff_tail));

	sb_1__1_ sb_7__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__64_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__66_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__63_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__57_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_54_ccff_tail),
		.chany_top_out(sb_1__1__57_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__57_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__57_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__57_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__57_ccff_tail));

	sb_1__1_ sb_7__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__65_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__67_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__64_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__58_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_75_ccff_tail),
		.chany_top_out(sb_1__1__58_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__58_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__58_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__58_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__58_ccff_tail));

	sb_1__1_ sb_7__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__66_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__68_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__65_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__59_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_56_ccff_tail),
		.chany_top_out(sb_1__1__59_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__59_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__59_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__59_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__59_ccff_tail));

	sb_1__1_ sb_7__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__67_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__69_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__66_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__60_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_77_ccff_tail),
		.chany_top_out(sb_1__1__60_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__60_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__60_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__60_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__60_ccff_tail));

	sb_1__1_ sb_7__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__68_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__70_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__67_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__61_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_58_ccff_tail),
		.chany_top_out(sb_1__1__61_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__61_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__61_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__61_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__61_ccff_tail));

	sb_1__1_ sb_7__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_1__1__69_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__1__71_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__68_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_78_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__62_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_79_ccff_tail),
		.chany_top_out(sb_1__1__62_chany_top_out[0:8]),
		.chanx_right_out(sb_1__1__62_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__1__62_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__1__62_chanx_left_out[0:8]),
		.ccff_tail(sb_1__1__62_ccff_tail));

	sb_1__10_ sb_1__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__1_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__0_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__10__0_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__0_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__0_ccff_tail));

	sb_1__10_ sb_2__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__2_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__1_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__10__1_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__1_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__1_ccff_tail));

	sb_1__10_ sb_3__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__3_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__2_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chanx_right_out(sb_1__10__2_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__2_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__2_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__2_ccff_tail));

	sb_1__10_ sb_4__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__4_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__3_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_4_ccff_tail),
		.chanx_right_out(sb_1__10__3_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__3_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__3_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__3_ccff_tail));

	sb_1__10_ sb_5__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__5_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__4_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_5_ccff_tail),
		.chanx_right_out(sb_1__10__4_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__4_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__4_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__4_ccff_tail));

	sb_1__10_ sb_6__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__6_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__59_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__5_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_6_ccff_tail),
		.chanx_right_out(sb_1__10__5_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__5_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__5_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__5_ccff_tail));

	sb_1__10_ sb_7__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_right_in(cbx_1__10__7_chanx_left_out[0:8]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__69_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_79_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__6_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_7_ccff_tail),
		.chanx_right_out(sb_1__10__6_chanx_right_out[0:8]),
		.chany_bottom_out(sb_1__10__6_chany_bottom_out[0:8]),
		.chanx_left_out(sb_1__10__6_chanx_left_out[0:8]),
		.ccff_tail(sb_1__10__6_ccff_tail));

	sb_8__0_ sb_8__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__0_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.ccff_head(grid_clb_60_ccff_tail),
		.chany_top_out(sb_8__0__0_chany_top_out[0:8]),
		.chanx_left_out(sb_8__0__0_chanx_left_out[0:8]),
		.ccff_tail(sb_8__0__0_ccff_tail));

	sb_8__1_ sb_8__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__1_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__0_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__63_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_70_ccff_tail),
		.chany_top_out(sb_8__1__0_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__0_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__0_ccff_tail));

	sb_8__1_ sb_8__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__2_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__1_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__64_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_62_ccff_tail),
		.chany_top_out(sb_8__1__1_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__1_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__1_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__1_ccff_tail));

	sb_8__1_ sb_8__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__3_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__2_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__65_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_72_ccff_tail),
		.chany_top_out(sb_8__1__2_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__2_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__2_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__2_ccff_tail));

	sb_8__1_ sb_8__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__4_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__3_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__66_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_64_ccff_tail),
		.chany_top_out(sb_8__1__3_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__3_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__3_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__3_ccff_tail));

	sb_8__1_ sb_8__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__5_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__4_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__67_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_74_ccff_tail),
		.chany_top_out(sb_8__1__4_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__4_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__4_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__4_ccff_tail));

	sb_8__1_ sb_8__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__6_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__5_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__68_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_66_ccff_tail),
		.chany_top_out(sb_8__1__5_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__5_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__5_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__5_ccff_tail));

	sb_8__1_ sb_8__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__7_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__6_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__69_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_76_ccff_tail),
		.chany_top_out(sb_8__1__6_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__6_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__6_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__6_ccff_tail));

	sb_8__1_ sb_8__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__8_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__7_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__70_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_78_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_68_ccff_tail),
		.chany_top_out(sb_8__1__7_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__7_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__7_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__7_ccff_tail));

	sb_8__1_ sb_8__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_top_in(cby_8__1__9_chany_bottom_out[0:8]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__8_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_78_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__71_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_79_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_78_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_78_ccff_tail),
		.chany_top_out(sb_8__1__8_chany_top_out[0:8]),
		.chany_bottom_out(sb_8__1__8_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__1__8_chanx_left_out[0:8]),
		.ccff_tail(sb_8__1__8_ccff_tail));

	sb_8__10_ sb_8__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(cby_8__1__9_chany_top_out[0:8]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_79_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__7_chanx_right_out[0:8]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_79_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_8__10__0_chany_bottom_out[0:8]),
		.chanx_left_out(sb_8__10__0_chanx_left_out[0:8]),
		.ccff_tail(sb_8__10__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__0__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__2_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__3_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__4_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__5_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__5_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:8]),
		.ccff_head(sb_1__0__6_ccff_tail),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__6_ccff_tail));

	cbx_1__0_ cbx_8__0_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__0__6_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__0__0_chanx_left_out[0:8]),
		.ccff_head(sb_8__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cbx_1__0__7_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_1__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__2_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_1__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__3_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_1__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__4_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_1__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__5_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__1_ cbx_1__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__6_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__6_ccff_tail));

	cbx_1__1_ cbx_1__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__7_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__7_ccff_tail));

	cbx_1__1_ cbx_1__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__1__8_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__8_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__9_ccff_tail),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__9_ccff_tail));

	cbx_1__1_ cbx_2__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__10_ccff_tail),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__10_ccff_tail));

	cbx_1__1_ cbx_2__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__2_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__11_ccff_tail),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__11_ccff_tail));

	cbx_1__1_ cbx_2__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__3_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__12_ccff_tail),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__12_ccff_tail));

	cbx_1__1_ cbx_2__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__4_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__13_ccff_tail),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__13_ccff_tail));

	cbx_1__1_ cbx_2__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__5_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__14_ccff_tail),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__14_ccff_tail));

	cbx_1__1_ cbx_2__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__6_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__15_ccff_tail),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__15_ccff_tail));

	cbx_1__1_ cbx_2__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__7_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__16_ccff_tail),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__16_ccff_tail));

	cbx_1__1_ cbx_2__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__8_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__17_ccff_tail),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__17_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__9_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__18_ccff_tail),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__18_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__10_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__19_ccff_tail),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__19_ccff_tail));

	cbx_1__1_ cbx_3__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__11_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__20_ccff_tail),
		.chanx_left_out(cbx_1__1__20_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__20_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__20_ccff_tail));

	cbx_1__1_ cbx_3__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__12_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__21_ccff_tail),
		.chanx_left_out(cbx_1__1__21_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__21_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__21_ccff_tail));

	cbx_1__1_ cbx_3__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__13_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__22_ccff_tail),
		.chanx_left_out(cbx_1__1__22_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__22_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__22_ccff_tail));

	cbx_1__1_ cbx_3__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__14_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__23_ccff_tail),
		.chanx_left_out(cbx_1__1__23_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__23_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__23_ccff_tail));

	cbx_1__1_ cbx_3__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__15_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__24_ccff_tail),
		.chanx_left_out(cbx_1__1__24_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__24_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__24_ccff_tail));

	cbx_1__1_ cbx_3__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__16_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__25_ccff_tail),
		.chanx_left_out(cbx_1__1__25_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__25_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__25_ccff_tail));

	cbx_1__1_ cbx_3__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__17_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__26_ccff_tail),
		.chanx_left_out(cbx_1__1__26_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__26_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__26_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__18_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__27_ccff_tail),
		.chanx_left_out(cbx_1__1__27_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__27_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__27_ccff_tail));

	cbx_1__1_ cbx_4__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__19_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__28_ccff_tail),
		.chanx_left_out(cbx_1__1__28_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__28_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__28_ccff_tail));

	cbx_1__1_ cbx_4__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__20_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__29_ccff_tail),
		.chanx_left_out(cbx_1__1__29_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__29_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__29_ccff_tail));

	cbx_1__1_ cbx_4__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__21_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__30_ccff_tail),
		.chanx_left_out(cbx_1__1__30_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__30_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__30_ccff_tail));

	cbx_1__1_ cbx_4__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__22_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__31_ccff_tail),
		.chanx_left_out(cbx_1__1__31_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__31_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__31_ccff_tail));

	cbx_1__1_ cbx_4__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__23_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__32_ccff_tail),
		.chanx_left_out(cbx_1__1__32_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__32_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__32_ccff_tail));

	cbx_1__1_ cbx_4__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__24_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__33_ccff_tail),
		.chanx_left_out(cbx_1__1__33_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__33_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__33_ccff_tail));

	cbx_1__1_ cbx_4__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__25_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__34_ccff_tail),
		.chanx_left_out(cbx_1__1__34_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__34_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__34_ccff_tail));

	cbx_1__1_ cbx_4__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__26_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__35_ccff_tail),
		.chanx_left_out(cbx_1__1__35_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__35_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__35_ccff_tail));

	cbx_1__1_ cbx_5__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__27_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__36_ccff_tail),
		.chanx_left_out(cbx_1__1__36_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__36_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__36_ccff_tail));

	cbx_1__1_ cbx_5__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__28_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__37_ccff_tail),
		.chanx_left_out(cbx_1__1__37_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__37_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__37_ccff_tail));

	cbx_1__1_ cbx_5__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__29_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__38_ccff_tail),
		.chanx_left_out(cbx_1__1__38_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__38_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__38_ccff_tail));

	cbx_1__1_ cbx_5__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__30_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__39_ccff_tail),
		.chanx_left_out(cbx_1__1__39_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__39_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__39_ccff_tail));

	cbx_1__1_ cbx_5__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__31_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__40_ccff_tail),
		.chanx_left_out(cbx_1__1__40_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__40_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__40_ccff_tail));

	cbx_1__1_ cbx_5__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__32_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__41_ccff_tail),
		.chanx_left_out(cbx_1__1__41_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__41_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__41_ccff_tail));

	cbx_1__1_ cbx_5__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__33_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__42_ccff_tail),
		.chanx_left_out(cbx_1__1__42_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__42_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__42_ccff_tail));

	cbx_1__1_ cbx_5__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__34_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__43_ccff_tail),
		.chanx_left_out(cbx_1__1__43_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__43_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__43_ccff_tail));

	cbx_1__1_ cbx_5__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__35_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__44_ccff_tail),
		.chanx_left_out(cbx_1__1__44_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__44_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__44_ccff_tail));

	cbx_1__1_ cbx_6__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__36_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__45_ccff_tail),
		.chanx_left_out(cbx_1__1__45_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__45_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__45_ccff_tail));

	cbx_1__1_ cbx_6__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__37_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__46_ccff_tail),
		.chanx_left_out(cbx_1__1__46_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__46_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__46_ccff_tail));

	cbx_1__1_ cbx_6__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__38_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__47_ccff_tail),
		.chanx_left_out(cbx_1__1__47_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__47_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__47_ccff_tail));

	cbx_1__1_ cbx_6__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__39_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__48_ccff_tail),
		.chanx_left_out(cbx_1__1__48_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__48_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__48_ccff_tail));

	cbx_1__1_ cbx_6__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__40_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__49_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__49_ccff_tail),
		.chanx_left_out(cbx_1__1__49_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__49_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__49_ccff_tail));

	cbx_1__1_ cbx_6__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__41_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__50_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__50_ccff_tail),
		.chanx_left_out(cbx_1__1__50_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__50_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__50_ccff_tail));

	cbx_1__1_ cbx_6__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__42_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__51_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__51_ccff_tail),
		.chanx_left_out(cbx_1__1__51_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__51_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__51_ccff_tail));

	cbx_1__1_ cbx_6__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__43_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__52_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__52_ccff_tail),
		.chanx_left_out(cbx_1__1__52_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__52_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__52_ccff_tail));

	cbx_1__1_ cbx_6__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__44_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__53_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__53_ccff_tail),
		.chanx_left_out(cbx_1__1__53_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__53_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__53_ccff_tail));

	cbx_1__1_ cbx_7__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__45_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__54_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__54_ccff_tail),
		.chanx_left_out(cbx_1__1__54_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__54_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__54_ccff_tail));

	cbx_1__1_ cbx_7__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__46_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__55_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__55_ccff_tail),
		.chanx_left_out(cbx_1__1__55_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__55_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__55_ccff_tail));

	cbx_1__1_ cbx_7__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__47_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__56_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__56_ccff_tail),
		.chanx_left_out(cbx_1__1__56_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__56_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__56_ccff_tail));

	cbx_1__1_ cbx_7__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__48_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__57_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__57_ccff_tail),
		.chanx_left_out(cbx_1__1__57_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__57_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__57_ccff_tail));

	cbx_1__1_ cbx_7__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__49_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__58_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__58_ccff_tail),
		.chanx_left_out(cbx_1__1__58_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__58_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__58_ccff_tail));

	cbx_1__1_ cbx_7__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__50_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__59_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__59_ccff_tail),
		.chanx_left_out(cbx_1__1__59_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__59_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__59_ccff_tail));

	cbx_1__1_ cbx_7__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__51_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__60_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__60_ccff_tail),
		.chanx_left_out(cbx_1__1__60_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__60_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__60_ccff_tail));

	cbx_1__1_ cbx_7__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__52_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__61_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__61_ccff_tail),
		.chanx_left_out(cbx_1__1__61_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__61_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__61_ccff_tail));

	cbx_1__1_ cbx_7__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__53_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__1__62_chanx_left_out[0:8]),
		.ccff_head(sb_1__1__62_ccff_tail),
		.chanx_left_out(cbx_1__1__62_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__62_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__62_ccff_tail));

	cbx_1__1_ cbx_8__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__54_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__0_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__63_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__63_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__63_ccff_tail));

	cbx_1__1_ cbx_8__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__55_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__1_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__64_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__64_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__64_ccff_tail));

	cbx_1__1_ cbx_8__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__56_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__2_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__65_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__65_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__65_ccff_tail));

	cbx_1__1_ cbx_8__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__57_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__3_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__66_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__66_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__66_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__66_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__66_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__66_ccff_tail));

	cbx_1__1_ cbx_8__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__58_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__4_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__67_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__67_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__67_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__67_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__67_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__67_ccff_tail));

	cbx_1__1_ cbx_8__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__59_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__5_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__68_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__68_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__68_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__68_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__68_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__68_ccff_tail));

	cbx_1__1_ cbx_8__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__60_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__6_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__69_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__69_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__69_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__69_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__69_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__69_ccff_tail));

	cbx_1__1_ cbx_8__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__61_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__7_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__7_ccff_tail),
		.chanx_left_out(cbx_1__1__70_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__70_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__70_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__70_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__70_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__70_ccff_tail));

	cbx_1__1_ cbx_8__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__1__62_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__1__8_chanx_left_out[0:8]),
		.ccff_head(sb_8__1__8_ccff_tail),
		.chanx_left_out(cbx_1__1__71_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__1__71_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__71_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__71_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__71_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__71_ccff_tail));

	cbx_1__10_ cbx_1__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_0__10__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__0_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__0_ccff_tail),
		.chanx_left_out(cbx_1__10__0_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__0_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__0_ccff_tail));

	cbx_1__10_ cbx_2__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__0_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__1_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__1_ccff_tail),
		.chanx_left_out(cbx_1__10__1_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__1_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__1_ccff_tail));

	cbx_1__10_ cbx_3__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__1_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__2_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__2_ccff_tail),
		.chanx_left_out(cbx_1__10__2_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__2_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__2_ccff_tail));

	cbx_1__10_ cbx_4__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__2_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__3_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__3_ccff_tail),
		.chanx_left_out(cbx_1__10__3_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__3_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__3_ccff_tail));

	cbx_1__10_ cbx_5__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__3_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__4_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__4_ccff_tail),
		.chanx_left_out(cbx_1__10__4_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__4_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__4_ccff_tail));

	cbx_1__10_ cbx_6__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__4_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__5_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__5_ccff_tail),
		.chanx_left_out(cbx_1__10__5_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__5_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__5_ccff_tail));

	cbx_1__10_ cbx_7__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__5_chanx_right_out[0:8]),
		.chanx_right_in(sb_1__10__6_chanx_left_out[0:8]),
		.ccff_head(sb_1__10__6_ccff_tail),
		.chanx_left_out(cbx_1__10__6_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__6_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__6_ccff_tail));

	cbx_1__10_ cbx_8__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chanx_left_in(sb_1__10__6_chanx_right_out[0:8]),
		.chanx_right_in(sb_8__10__0_chanx_left_out[0:8]),
		.ccff_head(sb_8__10__0_ccff_tail),
		.chanx_left_out(cbx_1__10__7_chanx_left_out[0:8]),
		.chanx_right_out(cbx_1__10__7_chanx_right_out[0:8]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__7_ccff_tail));

	cby_0__1_ cby_0__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:8]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__2_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__3_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__1_ cby_0__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__4_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__4_ccff_tail),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__5_ccff_tail));

	cby_0__1_ cby_0__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__5_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__5_ccff_tail),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__6_ccff_tail));

	cby_0__1_ cby_0__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__6_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__7_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__6_ccff_tail),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__7_ccff_tail));

	cby_0__1_ cby_0__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__7_chany_top_out[0:8]),
		.chany_top_in(sb_0__1__8_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__7_ccff_tail),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__8_ccff_tail));

	cby_0__1_ cby_0__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_0__1__8_chany_top_out[0:8]),
		.chany_top_in(sb_0__10__0_chany_bottom_out[0:8]),
		.ccff_head(sb_0__1__8_ccff_tail),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:8]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_tail(cby_0__1__9_ccff_tail));

	cby_1__1_ cby_1__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__2_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_1__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__3_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_1__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__4_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_1__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__5_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_1__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__6_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__6_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_1__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__7_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__7_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_1__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__8_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__8_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_2__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__1_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_2__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__9_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__9_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_1__1_ cby_2__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__10_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__10_ccff_tail),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__12_ccff_tail));

	cby_1__1_ cby_2__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__11_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__11_ccff_tail),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__13_ccff_tail));

	cby_1__1_ cby_2__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__12_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__12_ccff_tail),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__14_ccff_tail));

	cby_1__1_ cby_2__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__13_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__13_ccff_tail),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__15_ccff_tail));

	cby_1__1_ cby_2__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__14_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__14_ccff_tail),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__16_ccff_tail));

	cby_1__1_ cby_2__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__15_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__15_ccff_tail),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__17_ccff_tail));

	cby_1__1_ cby_2__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__16_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__16_ccff_tail),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__18_ccff_tail));

	cby_1__1_ cby_2__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__17_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__17_ccff_tail),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__19_ccff_tail));

	cby_1__1_ cby_3__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__2_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__20_ccff_tail));

	cby_1__1_ cby_3__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__18_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__18_ccff_tail),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__21_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__21_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__21_ccff_tail));

	cby_1__1_ cby_3__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__19_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__19_ccff_tail),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__22_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__22_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__22_ccff_tail));

	cby_1__1_ cby_3__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__20_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__20_ccff_tail),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__23_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__23_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__23_ccff_tail));

	cby_1__1_ cby_3__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__21_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__21_ccff_tail),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__24_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__24_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__24_ccff_tail));

	cby_1__1_ cby_3__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__22_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__22_ccff_tail),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__25_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__25_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__25_ccff_tail));

	cby_1__1_ cby_3__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__23_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__23_ccff_tail),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__26_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__26_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__26_ccff_tail));

	cby_1__1_ cby_3__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__24_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__24_ccff_tail),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__27_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__27_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__27_ccff_tail));

	cby_1__1_ cby_3__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__25_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__25_ccff_tail),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__28_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__28_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__28_ccff_tail));

	cby_1__1_ cby_3__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__26_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__2_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__26_ccff_tail),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__29_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__29_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__29_ccff_tail));

	cby_1__1_ cby_4__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__3_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__30_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__30_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__30_ccff_tail));

	cby_1__1_ cby_4__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__27_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__27_ccff_tail),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__31_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__31_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__31_ccff_tail));

	cby_1__1_ cby_4__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__28_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__28_ccff_tail),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__32_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__32_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__32_ccff_tail));

	cby_1__1_ cby_4__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__29_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__29_ccff_tail),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__33_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__33_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__33_ccff_tail));

	cby_1__1_ cby_4__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__30_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__30_ccff_tail),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__34_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__34_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__34_ccff_tail));

	cby_1__1_ cby_4__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__31_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__31_ccff_tail),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__35_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__35_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__35_ccff_tail));

	cby_1__1_ cby_4__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__32_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__32_ccff_tail),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__36_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__36_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__36_ccff_tail));

	cby_1__1_ cby_4__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__33_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__33_ccff_tail),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__37_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__37_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__37_ccff_tail));

	cby_1__1_ cby_4__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__34_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__34_ccff_tail),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__38_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__38_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__38_ccff_tail));

	cby_1__1_ cby_4__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__35_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__3_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__35_ccff_tail),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__39_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__39_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__39_ccff_tail));

	cby_1__1_ cby_5__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__4_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__40_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__40_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__40_ccff_tail));

	cby_1__1_ cby_5__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__36_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__36_ccff_tail),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__41_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__41_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__41_ccff_tail));

	cby_1__1_ cby_5__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__37_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__37_ccff_tail),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__42_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__42_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__42_ccff_tail));

	cby_1__1_ cby_5__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__38_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__38_ccff_tail),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__43_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__43_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__43_ccff_tail));

	cby_1__1_ cby_5__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__39_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__39_ccff_tail),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__44_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__44_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__44_ccff_tail));

	cby_1__1_ cby_5__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__40_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__40_ccff_tail),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__45_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__45_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__45_ccff_tail));

	cby_1__1_ cby_5__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__41_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__41_ccff_tail),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__46_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__46_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__46_ccff_tail));

	cby_1__1_ cby_5__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__42_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__42_ccff_tail),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__47_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__47_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__47_ccff_tail));

	cby_1__1_ cby_5__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__43_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__43_ccff_tail),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__48_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__48_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__48_ccff_tail));

	cby_1__1_ cby_5__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__44_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__4_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__44_ccff_tail),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__49_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__49_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__49_ccff_tail));

	cby_1__1_ cby_6__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__5_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__50_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__50_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__50_ccff_tail));

	cby_1__1_ cby_6__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__45_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__45_ccff_tail),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__51_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__51_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__51_ccff_tail));

	cby_1__1_ cby_6__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__46_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__46_ccff_tail),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__52_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__52_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__52_ccff_tail));

	cby_1__1_ cby_6__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__47_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__47_ccff_tail),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__53_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__53_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__53_ccff_tail));

	cby_1__1_ cby_6__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__48_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__49_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__48_ccff_tail),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__54_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__54_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__54_ccff_tail));

	cby_1__1_ cby_6__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__49_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__50_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__49_ccff_tail),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__55_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__55_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__55_ccff_tail));

	cby_1__1_ cby_6__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__50_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__51_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__50_ccff_tail),
		.chany_bottom_out(cby_1__1__56_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__56_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__56_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__56_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__56_ccff_tail));

	cby_1__1_ cby_6__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__51_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__52_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__51_ccff_tail),
		.chany_bottom_out(cby_1__1__57_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__57_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__57_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__57_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__57_ccff_tail));

	cby_1__1_ cby_6__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__52_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__53_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__52_ccff_tail),
		.chany_bottom_out(cby_1__1__58_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__58_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__58_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__58_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__58_ccff_tail));

	cby_1__1_ cby_6__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__53_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__5_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__53_ccff_tail),
		.chany_bottom_out(cby_1__1__59_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__59_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__59_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__59_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__59_ccff_tail));

	cby_1__1_ cby_7__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__0__6_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__54_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__6_ccff_tail),
		.chany_bottom_out(cby_1__1__60_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__60_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__60_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__60_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__60_ccff_tail));

	cby_1__1_ cby_7__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__54_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__55_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__54_ccff_tail),
		.chany_bottom_out(cby_1__1__61_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__61_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__61_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__61_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__61_ccff_tail));

	cby_1__1_ cby_7__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__55_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__56_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__55_ccff_tail),
		.chany_bottom_out(cby_1__1__62_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__62_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__62_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__62_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__62_ccff_tail));

	cby_1__1_ cby_7__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__56_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__57_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__56_ccff_tail),
		.chany_bottom_out(cby_1__1__63_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__63_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__63_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__63_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__63_ccff_tail));

	cby_1__1_ cby_7__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__57_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__58_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__57_ccff_tail),
		.chany_bottom_out(cby_1__1__64_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__64_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__64_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__64_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__64_ccff_tail));

	cby_1__1_ cby_7__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__58_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__59_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__58_ccff_tail),
		.chany_bottom_out(cby_1__1__65_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__65_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__65_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__65_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__65_ccff_tail));

	cby_1__1_ cby_7__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__59_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__60_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__59_ccff_tail),
		.chany_bottom_out(cby_1__1__66_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__66_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__66_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__66_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__66_ccff_tail));

	cby_1__1_ cby_7__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__60_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__61_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__60_ccff_tail),
		.chany_bottom_out(cby_1__1__67_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__67_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__67_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__67_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__67_ccff_tail));

	cby_1__1_ cby_7__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__61_chany_top_out[0:8]),
		.chany_top_in(sb_1__1__62_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__61_ccff_tail),
		.chany_bottom_out(cby_1__1__68_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__68_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__68_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__68_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__68_ccff_tail));

	cby_1__1_ cby_7__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_1__1__62_chany_top_out[0:8]),
		.chany_top_in(sb_1__10__6_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__62_ccff_tail),
		.chany_bottom_out(cby_1__1__69_chany_bottom_out[0:8]),
		.chany_top_out(cby_1__1__69_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__69_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__69_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__69_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__69_ccff_tail));

	cby_8__1_ cby_8__1_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__0__0_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__0__7_ccff_tail),
		.chany_bottom_out(cby_8__1__0_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__0_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__0_ccff_tail));

	cby_8__1_ cby_8__2_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__0_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__1_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__63_ccff_tail),
		.chany_bottom_out(cby_8__1__1_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__1_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__1_ccff_tail));

	cby_8__1_ cby_8__3_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__1_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__2_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__64_ccff_tail),
		.chany_bottom_out(cby_8__1__2_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__2_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__2_ccff_tail));

	cby_8__1_ cby_8__4_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__2_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__3_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__65_ccff_tail),
		.chany_bottom_out(cby_8__1__3_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__3_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__3_ccff_tail));

	cby_8__1_ cby_8__5_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__3_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__4_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__66_ccff_tail),
		.chany_bottom_out(cby_8__1__4_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__4_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__4_ccff_tail));

	cby_8__1_ cby_8__6_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__4_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__5_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__67_ccff_tail),
		.chany_bottom_out(cby_8__1__5_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__5_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__5_ccff_tail));

	cby_8__1_ cby_8__7_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__5_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__6_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__68_ccff_tail),
		.chany_bottom_out(cby_8__1__6_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__6_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__6_ccff_tail));

	cby_8__1_ cby_8__8_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__6_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__7_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__69_ccff_tail),
		.chany_bottom_out(cby_8__1__7_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__7_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__7_ccff_tail));

	cby_8__1_ cby_8__9_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__7_chany_top_out[0:8]),
		.chany_top_in(sb_8__1__8_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__70_ccff_tail),
		.chany_bottom_out(cby_8__1__8_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__8_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__8_ccff_tail));

	cby_8__1_ cby_8__10_ (
		`ifdef USE_POWER_PINS
  .vdd(vccd1),
  .vss(vssd1),
`endif
.prog_clk(prog_clk),

		.chany_bottom_in(sb_8__1__8_chany_top_out[0:8]),
		.chany_top_in(sb_8__10__0_chany_bottom_out[0:8]),
		.ccff_head(cbx_1__1__71_ccff_tail),
		.chany_bottom_out(cby_8__1__9_chany_bottom_out[0:8]),
		.chany_top_out(cby_8__1__9_chany_top_out[0:8]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_8__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_8__1__9_ccff_tail));


// ----- END Verilog module for fpga_top -----






endmodule	// user_project_wrapper

`default_nettype wire
