// This is the unpowered netlist.
module grid_clb (bottom_width_0_height_0_subtile_0__pin_I_2_,
    bottom_width_0_height_0_subtile_0__pin_I_6_,
    bottom_width_0_height_0_subtile_0__pin_O_0_,
    bottom_width_0_height_0_subtile_0__pin_clk_0_,
    ccff_head,
    ccff_tail,
    clk,
    left_width_0_height_0_subtile_0__pin_I_3_,
    left_width_0_height_0_subtile_0__pin_I_7_,
    left_width_0_height_0_subtile_0__pin_O_1_,
    prog_clk,
    reset,
    right_width_0_height_0_subtile_0__pin_I_1_,
    right_width_0_height_0_subtile_0__pin_I_5_,
    right_width_0_height_0_subtile_0__pin_I_9_,
    right_width_0_height_0_subtile_0__pin_O_3_,
    set,
    top_width_0_height_0_subtile_0__pin_I_0_,
    top_width_0_height_0_subtile_0__pin_I_4_,
    top_width_0_height_0_subtile_0__pin_I_8_,
    top_width_0_height_0_subtile_0__pin_O_2_);
 input bottom_width_0_height_0_subtile_0__pin_I_2_;
 input bottom_width_0_height_0_subtile_0__pin_I_6_;
 output bottom_width_0_height_0_subtile_0__pin_O_0_;
 input bottom_width_0_height_0_subtile_0__pin_clk_0_;
 input ccff_head;
 output ccff_tail;
 input clk;
 input left_width_0_height_0_subtile_0__pin_I_3_;
 input left_width_0_height_0_subtile_0__pin_I_7_;
 output left_width_0_height_0_subtile_0__pin_O_1_;
 input prog_clk;
 input reset;
 input right_width_0_height_0_subtile_0__pin_I_1_;
 input right_width_0_height_0_subtile_0__pin_I_5_;
 input right_width_0_height_0_subtile_0__pin_I_9_;
 output right_width_0_height_0_subtile_0__pin_O_3_;
 input set;
 input top_width_0_height_0_subtile_0__pin_I_0_;
 input top_width_0_height_0_subtile_0__pin_I_4_;
 input top_width_0_height_0_subtile_0__pin_I_8_;
 output top_width_0_height_0_subtile_0__pin_O_2_;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire clknet_0_prog_clk;
 wire clknet_4_0_0_prog_clk;
 wire clknet_4_10_0_prog_clk;
 wire clknet_4_11_0_prog_clk;
 wire clknet_4_12_0_prog_clk;
 wire clknet_4_13_0_prog_clk;
 wire clknet_4_14_0_prog_clk;
 wire clknet_4_15_0_prog_clk;
 wire clknet_4_1_0_prog_clk;
 wire clknet_4_2_0_prog_clk;
 wire clknet_4_3_0_prog_clk;
 wire clknet_4_4_0_prog_clk;
 wire clknet_4_5_0_prog_clk;
 wire clknet_4_6_0_prog_clk;
 wire clknet_4_7_0_prog_clk;
 wire clknet_4_8_0_prog_clk;
 wire clknet_4_9_0_prog_clk;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ;
 wire \logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out ;
 wire \logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(right_width_0_height_0_subtile_0__pin_I_5_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_60 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__clkinv_4 _0928_ (.A(net7),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _0929_ (.A(_0009_),
    .B(net11),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _0930_ (.A(_0009_),
    .B(net11),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0931_ (.A(net7),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_1 _0932_ (.A(_0009_),
    .B(net11),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0933_ (.A(net7),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _0934_ (.A(_0009_),
    .B(net11),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0935_ (.A(net7),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0936_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .Y(_0890_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_1 _0938_ (.A(_0276_),
    .X(_0891_));
 sky130_fd_sc_hd__inv_2 _0939_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0941_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0335_));
 sky130_fd_sc_hd__buf_6 _0942_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0277_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(_0277_),
    .Y(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0944_ (.A(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_1 _0945_ (.A(_0278_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_1 _0946_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0279_),
    .X(_0904_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(_0277_),
    .Y(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0277_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _0950_ (.A(_0280_),
    .X(_0899_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _0952_ (.A(_0281_),
    .X(_0906_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(_0277_),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0282_));
 sky130_fd_sc_hd__buf_1 _0956_ (.A(_0282_),
    .X(_0898_));
 sky130_fd_sc_hd__buf_1 _0957_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0283_));
 sky130_fd_sc_hd__buf_1 _0958_ (.A(_0283_),
    .X(_0903_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(_0277_),
    .Y(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0284_));
 sky130_fd_sc_hd__buf_1 _0961_ (.A(_0284_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _0963_ (.A(_0285_),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0965_ (.A(_0286_),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0967_ (.A(_0287_),
    .X(_0701_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .Y(_0687_));
 sky130_fd_sc_hd__buf_6 _0969_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0970_ (.A(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0971_ (.A(_0289_),
    .X(_0697_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(_0288_),
    .Y(_0683_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .Y(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0975_ (.A(_0290_),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(_0288_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0291_),
    .X(_0696_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(_0288_),
    .Y(_0682_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .Y(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0288_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0981_ (.A(_0292_),
    .X(_0695_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(_0288_),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .Y(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _0984_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0293_),
    .X(_0702_));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(_0294_),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(_0295_),
    .X(_0694_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0288_),
    .Y(_0680_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .Y(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(_0296_),
    .X(_0693_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(_0288_),
    .Y(_0679_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .Y(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(_0297_),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(_0298_),
    .X(_0692_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(_0288_),
    .Y(_0678_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .Y(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0299_),
    .X(_0691_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(_0288_),
    .Y(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(_0300_),
    .X(_0907_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(_0277_),
    .Y(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(_0301_),
    .X(_0896_));
 sky130_fd_sc_hd__buf_1 _1012_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0302_));
 sky130_fd_sc_hd__buf_1 _1013_ (.A(_0302_),
    .X(_0902_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(_0277_),
    .Y(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _1016_ (.A(_0303_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .X(_0304_));
 sky130_fd_sc_hd__buf_1 _1018_ (.A(_0304_),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(_0305_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(_0306_),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .Y(_0715_));
 sky130_fd_sc_hd__buf_6 _1024_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _1026_ (.A(_0308_),
    .X(_0725_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(_0307_),
    .Y(_0711_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .Y(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(_0309_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0307_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(_0310_),
    .X(_0724_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(_0307_),
    .Y(_0710_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .Y(_0714_));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(_0307_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0311_),
    .X(_0723_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(_0307_),
    .Y(_0709_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .Y(_0718_));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0312_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _1042_ (.A(_0313_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_1 _1043_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _1044_ (.A(_0314_),
    .X(_0722_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0307_),
    .Y(_0708_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .Y(_0713_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _1048_ (.A(_0315_),
    .X(_0721_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0307_),
    .Y(_0707_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .Y(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _1052_ (.A(_0316_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _1054_ (.A(_0317_),
    .X(_0720_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0307_),
    .Y(_0706_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .Y(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _1057_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _1058_ (.A(_0318_),
    .X(_0719_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0307_),
    .Y(_0705_));
 sky130_fd_sc_hd__clkbuf_1 _1060_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0319_),
    .X(_0905_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0277_),
    .Y(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _1064_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0320_),
    .X(_0894_));
 sky130_fd_sc_hd__clkbuf_1 _1066_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .X(_0321_));
 sky130_fd_sc_hd__buf_1 _1067_ (.A(_0321_),
    .X(_0760_));
 sky130_fd_sc_hd__clkbuf_1 _1068_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _1069_ (.A(_0322_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _1071_ (.A(_0323_),
    .X(_0757_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .Y(_0743_));
 sky130_fd_sc_hd__buf_6 _1073_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(_0012_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(_0013_),
    .X(_0753_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0012_),
    .Y(_0739_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .Y(_0745_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_1 _1079_ (.A(_0014_),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_1 _1080_ (.A(_0012_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_1 _1081_ (.A(_0015_),
    .X(_0752_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(_0012_),
    .Y(_0738_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .Y(_0742_));
 sky130_fd_sc_hd__clkbuf_1 _1084_ (.A(_0012_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_1 _1085_ (.A(_0016_),
    .X(_0751_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(_0012_),
    .Y(_0737_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .Y(_0746_));
 sky130_fd_sc_hd__clkbuf_1 _1088_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0017_),
    .X(_0758_));
 sky130_fd_sc_hd__clkbuf_1 _1090_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_1 _1091_ (.A(_0018_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _1092_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_1 _1093_ (.A(_0019_),
    .X(_0750_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(_0012_),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .Y(_0741_));
 sky130_fd_sc_hd__clkbuf_1 _1096_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_1 _1097_ (.A(_0020_),
    .X(_0749_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(_0012_),
    .Y(_0735_));
 sky130_fd_sc_hd__inv_2 _1099_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .Y(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _1100_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_1 _1101_ (.A(_0021_),
    .X(_0754_));
 sky130_fd_sc_hd__clkbuf_1 _1102_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_1 _1103_ (.A(_0022_),
    .X(_0748_));
 sky130_fd_sc_hd__inv_2 _1104_ (.A(_0012_),
    .Y(_0734_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .Y(_0740_));
 sky130_fd_sc_hd__clkbuf_1 _1106_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_1 _1107_ (.A(_0023_),
    .X(_0747_));
 sky130_fd_sc_hd__inv_2 _1108_ (.A(_0012_),
    .Y(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _1109_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_1 _1110_ (.A(_0024_),
    .X(_0901_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(_0277_),
    .Y(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _1112_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .X(_0025_));
 sky130_fd_sc_hd__buf_1 _1113_ (.A(_0025_),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_1 _1115_ (.A(_0026_),
    .X(_0787_));
 sky130_fd_sc_hd__clkbuf_1 _1116_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_1 _1117_ (.A(_0027_),
    .X(_0785_));
 sky130_fd_sc_hd__inv_2 _1118_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .Y(_0771_));
 sky130_fd_sc_hd__buf_6 _1119_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_1 _1120_ (.A(_0028_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_1 _1121_ (.A(_0029_),
    .X(_0781_));
 sky130_fd_sc_hd__inv_2 _1122_ (.A(_0028_),
    .Y(_0767_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .Y(_0773_));
 sky130_fd_sc_hd__clkbuf_1 _1124_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_1 _1125_ (.A(_0030_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_1 _1126_ (.A(_0028_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_1 _1127_ (.A(_0031_),
    .X(_0780_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .Y(_0856_));
 sky130_fd_sc_hd__clkbuf_1 _1129_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(_0032_));
 sky130_fd_sc_hd__clkbuf_1 _1130_ (.A(_0032_),
    .X(_0857_));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .Y(_0888_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0885_));
 sky130_fd_sc_hd__buf_6 _1134_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(_0033_),
    .Y(_0881_));
 sky130_fd_sc_hd__clkbuf_1 _1136_ (.A(_0033_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0034_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_1 _1138_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_1 _1139_ (.A(_0035_),
    .X(_0870_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(_0033_),
    .Y(_0880_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0033_),
    .X(_0036_));
 sky130_fd_sc_hd__clkbuf_1 _1142_ (.A(_0036_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _1143_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_1 _1144_ (.A(_0037_),
    .X(_0872_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0884_));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(_0033_),
    .Y(_0879_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_1 _1148_ (.A(_0038_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_1 _1150_ (.A(_0039_),
    .X(_0869_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(_0033_),
    .Y(_0878_));
 sky130_fd_sc_hd__clkbuf_1 _1152_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0040_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0040_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_1 _1154_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_1 _1155_ (.A(_0041_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_1 _1156_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_1 _1157_ (.A(_0042_),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_1 _1158_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_1 _1159_ (.A(_0043_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .Y(_0575_));
 sky130_fd_sc_hd__buf_6 _1161_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_1 _1162_ (.A(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_1 _1163_ (.A(_0045_),
    .X(_0585_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(_0044_),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .Y(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1166_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_1 _1167_ (.A(_0046_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_1 _1168_ (.A(_0044_),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0047_),
    .X(_0584_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(_0044_),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .Y(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _1172_ (.A(_0044_),
    .X(_0048_));
 sky130_fd_sc_hd__clkbuf_1 _1173_ (.A(_0048_),
    .X(_0583_));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(_0044_),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_2 _1175_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .Y(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _1176_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_1 _1177_ (.A(_0049_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_1 _1178_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_1 _1179_ (.A(_0050_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _1180_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0051_),
    .X(_0582_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(_0044_),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .Y(_0573_));
 sky130_fd_sc_hd__clkbuf_1 _1184_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_1 _1185_ (.A(_0052_),
    .X(_0581_));
 sky130_fd_sc_hd__inv_2 _1186_ (.A(_0044_),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_2 _1187_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .Y(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _1188_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0053_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_1 _1190_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0054_),
    .X(_0580_));
 sky130_fd_sc_hd__inv_2 _1192_ (.A(_0044_),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .Y(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _1194_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_1 _1195_ (.A(_0055_),
    .X(_0579_));
 sky130_fd_sc_hd__inv_2 _1196_ (.A(_0044_),
    .Y(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1197_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .X(_0056_));
 sky130_fd_sc_hd__clkbuf_1 _1198_ (.A(_0056_),
    .X(_0873_));
 sky130_fd_sc_hd__inv_2 _1199_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0886_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(_0033_),
    .Y(_0877_));
 sky130_fd_sc_hd__clkbuf_1 _1202_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_1 _1203_ (.A(_0057_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _1204_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0058_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0058_),
    .X(_0868_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(_0033_),
    .Y(_0876_));
 sky130_fd_sc_hd__clkbuf_1 _1207_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_1 _1208_ (.A(_0059_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_1 _1209_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .X(_0060_));
 sky130_fd_sc_hd__buf_1 _1210_ (.A(_0060_),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_1 _1211_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_1 _1212_ (.A(_0061_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_1 _1213_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .X(_0062_));
 sky130_fd_sc_hd__clkbuf_1 _1214_ (.A(_0062_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _1215_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .Y(_0603_));
 sky130_fd_sc_hd__buf_6 _1216_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_1 _1217_ (.A(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_1 _1218_ (.A(_0064_),
    .X(_0613_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(_0063_),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _1220_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .Y(_0605_));
 sky130_fd_sc_hd__clkbuf_1 _1221_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_1 _1222_ (.A(_0065_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_1 _1223_ (.A(_0063_),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_1 _1224_ (.A(_0066_),
    .X(_0612_));
 sky130_fd_sc_hd__inv_2 _1225_ (.A(_0063_),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _1226_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .Y(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _1227_ (.A(_0063_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_1 _1228_ (.A(_0067_),
    .X(_0611_));
 sky130_fd_sc_hd__inv_2 _1229_ (.A(_0063_),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _1230_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .Y(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _1231_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_1 _1232_ (.A(_0068_),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_1 _1233_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_1 _1234_ (.A(_0069_),
    .X(_0615_));
 sky130_fd_sc_hd__clkbuf_1 _1235_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_1 _1236_ (.A(_0070_),
    .X(_0610_));
 sky130_fd_sc_hd__inv_2 _1237_ (.A(_0063_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _1238_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .Y(_0601_));
 sky130_fd_sc_hd__clkbuf_1 _1239_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_1 _1240_ (.A(_0071_),
    .X(_0609_));
 sky130_fd_sc_hd__inv_2 _1241_ (.A(_0063_),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _1242_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .Y(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _1243_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_1 _1244_ (.A(_0072_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _1245_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_1 _1246_ (.A(_0073_),
    .X(_0608_));
 sky130_fd_sc_hd__inv_2 _1247_ (.A(_0063_),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _1248_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .Y(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _1249_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_1 _1250_ (.A(_0074_),
    .X(_0607_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(_0063_),
    .Y(_0593_));
 sky130_fd_sc_hd__clkbuf_1 _1252_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_1 _1253_ (.A(_0075_),
    .X(_0871_));
 sky130_fd_sc_hd__inv_2 _1254_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(_0033_),
    .Y(_0875_));
 sky130_fd_sc_hd__clkbuf_1 _1256_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_1 _1257_ (.A(_0076_),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_1 _1258_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .X(_0077_));
 sky130_fd_sc_hd__buf_1 _1259_ (.A(_0077_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_1 _1260_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _1261_ (.A(_0078_),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_1 _1262_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(_0079_),
    .X(_0645_));
 sky130_fd_sc_hd__inv_2 _1264_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .Y(_0631_));
 sky130_fd_sc_hd__buf_6 _1265_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _1266_ (.A(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _1267_ (.A(_0081_),
    .X(_0641_));
 sky130_fd_sc_hd__inv_2 _1268_ (.A(_0080_),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _1269_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .Y(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1270_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _1271_ (.A(_0082_),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_1 _1272_ (.A(_0080_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _1273_ (.A(_0083_),
    .X(_0640_));
 sky130_fd_sc_hd__inv_2 _1274_ (.A(_0080_),
    .Y(_0626_));
 sky130_fd_sc_hd__inv_2 _1275_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .Y(_0630_));
 sky130_fd_sc_hd__clkbuf_1 _1276_ (.A(_0080_),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _1277_ (.A(_0084_),
    .X(_0639_));
 sky130_fd_sc_hd__inv_2 _1278_ (.A(_0080_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .Y(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _1280_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _1281_ (.A(_0085_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _1282_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _1283_ (.A(_0086_),
    .X(_0643_));
 sky130_fd_sc_hd__clkbuf_1 _1284_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _1285_ (.A(_0087_),
    .X(_0638_));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(_0080_),
    .Y(_0624_));
 sky130_fd_sc_hd__inv_2 _1287_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .Y(_0629_));
 sky130_fd_sc_hd__clkbuf_1 _1288_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _1289_ (.A(_0088_),
    .X(_0637_));
 sky130_fd_sc_hd__inv_2 _1290_ (.A(_0080_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _1291_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .Y(_0632_));
 sky130_fd_sc_hd__clkbuf_1 _1292_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _1293_ (.A(_0089_),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_1 _1294_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _1295_ (.A(_0090_),
    .X(_0636_));
 sky130_fd_sc_hd__inv_2 _1296_ (.A(_0080_),
    .Y(_0622_));
 sky130_fd_sc_hd__inv_2 _1297_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .Y(_0628_));
 sky130_fd_sc_hd__clkbuf_1 _1298_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _1299_ (.A(_0091_),
    .X(_0635_));
 sky130_fd_sc_hd__inv_2 _1300_ (.A(_0080_),
    .Y(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _1301_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _1302_ (.A(_0092_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(_0033_),
    .Y(_0874_));
 sky130_fd_sc_hd__clkbuf_1 _1304_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__buf_1 _1305_ (.A(_0093_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_1 _1306_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _1307_ (.A(_0094_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _1308_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _1309_ (.A(_0095_),
    .X(_0673_));
 sky130_fd_sc_hd__inv_2 _1310_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .Y(_0659_));
 sky130_fd_sc_hd__buf_6 _1311_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _1312_ (.A(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(_0097_),
    .X(_0669_));
 sky130_fd_sc_hd__inv_2 _1314_ (.A(_0096_),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_2 _1315_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .Y(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _1316_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _1317_ (.A(_0098_),
    .X(_0823_));
 sky130_fd_sc_hd__inv_2 _1318_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_2 _1319_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0851_));
 sky130_fd_sc_hd__buf_6 _1321_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0099_));
 sky130_fd_sc_hd__inv_2 _1322_ (.A(_0099_),
    .Y(_0847_));
 sky130_fd_sc_hd__clkbuf_1 _1323_ (.A(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _1324_ (.A(_0100_),
    .X(_0832_));
 sky130_fd_sc_hd__clkbuf_1 _1325_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _1326_ (.A(_0101_),
    .X(_0836_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(_0099_),
    .Y(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _1328_ (.A(_0099_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _1329_ (.A(_0102_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _1330_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _1331_ (.A(_0103_),
    .X(_0838_));
 sky130_fd_sc_hd__inv_2 _1332_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _1333_ (.A(_0099_),
    .Y(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _1334_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _1335_ (.A(_0104_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_1 _1336_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_1 _1337_ (.A(_0105_),
    .X(_0835_));
 sky130_fd_sc_hd__inv_2 _1338_ (.A(_0099_),
    .Y(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _1339_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _1340_ (.A(_0106_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_1 _1341_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _1342_ (.A(_0107_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _1344_ (.A(_0108_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _1345_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _1346_ (.A(_0109_),
    .X(_0477_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .Y(_0463_));
 sky130_fd_sc_hd__buf_6 _1348_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _1349_ (.A(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _1350_ (.A(_0111_),
    .X(_0473_));
 sky130_fd_sc_hd__inv_2 _1351_ (.A(_0110_),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .Y(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _1353_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _1354_ (.A(_0112_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _1355_ (.A(_0110_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _1356_ (.A(_0113_),
    .X(_0472_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(_0110_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .Y(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _1359_ (.A(_0110_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _1360_ (.A(_0114_),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(_0110_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _1362_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .Y(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _1363_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _1364_ (.A(_0115_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _1365_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _1366_ (.A(_0116_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1367_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _1368_ (.A(_0117_),
    .X(_0470_));
 sky130_fd_sc_hd__inv_2 _1369_ (.A(_0110_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _1370_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .Y(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _1371_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(_0118_),
    .X(_0469_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(_0110_),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .Y(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _1375_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(_0119_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _1377_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _1378_ (.A(_0120_),
    .X(_0468_));
 sky130_fd_sc_hd__inv_2 _1379_ (.A(_0110_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .Y(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _1381_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _1382_ (.A(_0121_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _1383_ (.A(_0110_),
    .Y(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _1384_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _1385_ (.A(_0122_),
    .X(_0839_));
 sky130_fd_sc_hd__inv_2 _1386_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _1387_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0849_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(_0099_),
    .Y(_0843_));
 sky130_fd_sc_hd__clkbuf_1 _1389_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _1390_ (.A(_0123_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _1391_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _1392_ (.A(_0124_),
    .X(_0834_));
 sky130_fd_sc_hd__inv_2 _1393_ (.A(_0099_),
    .Y(_0842_));
 sky130_fd_sc_hd__clkbuf_1 _1394_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _1395_ (.A(_0125_),
    .X(_0827_));
 sky130_fd_sc_hd__clkbuf_1 _1396_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .X(_0126_));
 sky130_fd_sc_hd__buf_1 _1397_ (.A(_0126_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1398_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _1399_ (.A(_0127_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1400_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _1401_ (.A(_0128_),
    .X(_0505_));
 sky130_fd_sc_hd__inv_2 _1402_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .Y(_0491_));
 sky130_fd_sc_hd__buf_6 _1403_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _1404_ (.A(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _1405_ (.A(_0130_),
    .X(_0501_));
 sky130_fd_sc_hd__inv_2 _1406_ (.A(_0129_),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_2 _1407_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .Y(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _1408_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _1409_ (.A(_0131_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _1410_ (.A(_0129_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _1411_ (.A(_0132_),
    .X(_0500_));
 sky130_fd_sc_hd__inv_2 _1412_ (.A(_0129_),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _1413_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .Y(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _1414_ (.A(_0129_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _1415_ (.A(_0133_),
    .X(_0499_));
 sky130_fd_sc_hd__inv_2 _1416_ (.A(_0129_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _1417_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .Y(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _1418_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _1419_ (.A(_0134_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _1420_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _1421_ (.A(_0135_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _1422_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1423_ (.A(_0136_),
    .X(_0498_));
 sky130_fd_sc_hd__inv_2 _1424_ (.A(_0129_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _1425_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .Y(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _1426_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _1427_ (.A(_0137_),
    .X(_0497_));
 sky130_fd_sc_hd__inv_2 _1428_ (.A(_0129_),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _1429_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .Y(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _1430_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1431_ (.A(_0138_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1432_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _1433_ (.A(_0139_),
    .X(_0496_));
 sky130_fd_sc_hd__inv_2 _1434_ (.A(_0129_),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _1435_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .Y(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _1436_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _1437_ (.A(_0140_),
    .X(_0495_));
 sky130_fd_sc_hd__inv_2 _1438_ (.A(_0129_),
    .Y(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _1439_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _1440_ (.A(_0141_),
    .X(_0837_));
 sky130_fd_sc_hd__inv_2 _1441_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0848_));
 sky130_fd_sc_hd__inv_2 _1442_ (.A(_0099_),
    .Y(_0841_));
 sky130_fd_sc_hd__clkbuf_1 _1443_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _1444_ (.A(_0142_),
    .X(_0826_));
 sky130_fd_sc_hd__clkbuf_1 _1445_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__buf_1 _1446_ (.A(_0143_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1447_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _1448_ (.A(_0144_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1449_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(_0145_),
    .X(_0533_));
 sky130_fd_sc_hd__inv_2 _1451_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .Y(_0519_));
 sky130_fd_sc_hd__buf_6 _1452_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _1453_ (.A(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _1454_ (.A(_0147_),
    .X(_0529_));
 sky130_fd_sc_hd__inv_2 _1455_ (.A(_0146_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _1456_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .Y(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _1457_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _1458_ (.A(_0148_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1459_ (.A(_0146_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _1460_ (.A(_0149_),
    .X(_0528_));
 sky130_fd_sc_hd__inv_2 _1461_ (.A(_0146_),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _1462_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .Y(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1463_ (.A(_0146_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _1464_ (.A(_0150_),
    .X(_0527_));
 sky130_fd_sc_hd__inv_2 _1465_ (.A(_0146_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _1466_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .Y(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _1467_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0151_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1469_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _1470_ (.A(_0152_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _1471_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _1472_ (.A(_0153_),
    .X(_0526_));
 sky130_fd_sc_hd__inv_2 _1473_ (.A(_0146_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _1474_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .Y(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1475_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _1476_ (.A(_0154_),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _1477_ (.A(_0146_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _1478_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .Y(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _1479_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _1480_ (.A(_0155_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1481_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _1482_ (.A(_0156_),
    .X(_0524_));
 sky130_fd_sc_hd__inv_2 _1483_ (.A(_0146_),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _1484_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .Y(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1485_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _1486_ (.A(_0157_),
    .X(_0523_));
 sky130_fd_sc_hd__inv_2 _1487_ (.A(_0146_),
    .Y(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1488_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _1489_ (.A(_0158_),
    .X(_0833_));
 sky130_fd_sc_hd__inv_2 _1490_ (.A(_0099_),
    .Y(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _1491_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__buf_1 _1492_ (.A(_0159_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _1493_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _1494_ (.A(_0160_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _1495_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0161_),
    .X(_0561_));
 sky130_fd_sc_hd__inv_2 _1497_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .Y(_0547_));
 sky130_fd_sc_hd__buf_6 _1498_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _1499_ (.A(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _1500_ (.A(_0163_),
    .X(_0557_));
 sky130_fd_sc_hd__inv_2 _1501_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _1502_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .Y(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _1503_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _1504_ (.A(_0164_),
    .X(_0789_));
 sky130_fd_sc_hd__inv_2 _1505_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_2 _1506_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _1507_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0817_));
 sky130_fd_sc_hd__buf_6 _1508_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0165_));
 sky130_fd_sc_hd__inv_2 _1509_ (.A(_0165_),
    .Y(_0813_));
 sky130_fd_sc_hd__clkbuf_1 _1510_ (.A(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _1511_ (.A(_0166_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_1 _1512_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _1513_ (.A(_0167_),
    .X(_0802_));
 sky130_fd_sc_hd__inv_2 _1514_ (.A(_0165_),
    .Y(_0812_));
 sky130_fd_sc_hd__clkbuf_1 _1515_ (.A(_0165_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _1516_ (.A(_0168_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_1 _1517_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_0169_),
    .X(_0804_));
 sky130_fd_sc_hd__inv_2 _1519_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _1520_ (.A(_0165_),
    .Y(_0811_));
 sky130_fd_sc_hd__clkbuf_1 _1521_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _1522_ (.A(_0170_),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_1 _1523_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _1524_ (.A(_0171_),
    .X(_0801_));
 sky130_fd_sc_hd__inv_2 _1525_ (.A(_0165_),
    .Y(_0810_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _1527_ (.A(_0172_),
    .X(_0795_));
 sky130_fd_sc_hd__clkbuf_1 _1528_ (.A(net16),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _1529_ (.A(_0173_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _1530_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _1531_ (.A(_0174_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _1533_ (.A(_0175_),
    .X(_0365_));
 sky130_fd_sc_hd__inv_2 _1534_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .Y(_0351_));
 sky130_fd_sc_hd__buf_6 _1535_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _1536_ (.A(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _1537_ (.A(_0177_),
    .X(_0361_));
 sky130_fd_sc_hd__inv_2 _1538_ (.A(_0176_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _1539_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .Y(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _1540_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0178_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _1542_ (.A(_0176_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _1543_ (.A(_0179_),
    .X(_0360_));
 sky130_fd_sc_hd__inv_2 _1544_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0176_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _1546_ (.A(_0180_),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _1547_ (.A(net16),
    .Y(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _1548_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _1549_ (.A(_0181_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _1550_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_1 _1551_ (.A(_0182_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _1552_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _1553_ (.A(_0183_),
    .X(_0358_));
 sky130_fd_sc_hd__inv_2 _1554_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .Y(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _1555_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _1556_ (.A(_0184_),
    .X(_0357_));
 sky130_fd_sc_hd__inv_2 _1557_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .Y(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _1558_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _1559_ (.A(_0185_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _1560_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _1561_ (.A(_0186_),
    .X(_0356_));
 sky130_fd_sc_hd__inv_2 _1562_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .Y(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _1563_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _1564_ (.A(_0187_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _1565_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1566_ (.A(_0188_),
    .X(_0805_));
 sky130_fd_sc_hd__inv_2 _1567_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _1568_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _1569_ (.A(_0165_),
    .Y(_0809_));
 sky130_fd_sc_hd__clkbuf_1 _1570_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1571_ (.A(_0189_),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_1 _1572_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _1573_ (.A(_0190_),
    .X(_0800_));
 sky130_fd_sc_hd__inv_2 _1574_ (.A(_0165_),
    .Y(_0808_));
 sky130_fd_sc_hd__clkbuf_1 _1575_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1576_ (.A(_0191_),
    .X(_0793_));
 sky130_fd_sc_hd__clkbuf_1 _1577_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .X(_0192_));
 sky130_fd_sc_hd__buf_1 _1578_ (.A(_0192_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1579_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _1580_ (.A(_0193_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1581_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _1582_ (.A(_0194_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _1583_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .Y(_0379_));
 sky130_fd_sc_hd__buf_6 _1584_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1585_ (.A(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _1586_ (.A(_0196_),
    .X(_0389_));
 sky130_fd_sc_hd__inv_2 _1587_ (.A(_0195_),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _1588_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .Y(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _1589_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1590_ (.A(_0197_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _1591_ (.A(_0195_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _1592_ (.A(_0198_),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _1593_ (.A(_0195_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _1594_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .Y(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _1595_ (.A(_0195_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_0199_),
    .X(_0387_));
 sky130_fd_sc_hd__inv_2 _1597_ (.A(_0195_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _1598_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .Y(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _1599_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _1600_ (.A(_0200_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _1601_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _1602_ (.A(_0201_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _1603_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _1604_ (.A(_0202_),
    .X(_0386_));
 sky130_fd_sc_hd__inv_2 _1605_ (.A(_0195_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _1606_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .Y(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _1607_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _1608_ (.A(_0203_),
    .X(_0385_));
 sky130_fd_sc_hd__inv_2 _1609_ (.A(_0195_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _1610_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .Y(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _1611_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _1612_ (.A(_0204_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _1613_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _1614_ (.A(_0205_),
    .X(_0384_));
 sky130_fd_sc_hd__inv_2 _1615_ (.A(_0195_),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _1616_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .Y(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _1617_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1618_ (.A(_0206_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _1619_ (.A(_0195_),
    .Y(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _1620_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _1621_ (.A(_0207_),
    .X(_0803_));
 sky130_fd_sc_hd__inv_2 _1622_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _1623_ (.A(_0165_),
    .Y(_0807_));
 sky130_fd_sc_hd__clkbuf_1 _1624_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _1625_ (.A(_0208_),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_1 _1626_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__buf_1 _1627_ (.A(_0209_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _1628_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _1629_ (.A(_0210_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _1630_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _1631_ (.A(_0211_),
    .X(_0421_));
 sky130_fd_sc_hd__inv_2 _1632_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .Y(_0407_));
 sky130_fd_sc_hd__buf_6 _1633_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1634_ (.A(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_1 _1635_ (.A(_0213_),
    .X(_0417_));
 sky130_fd_sc_hd__inv_2 _1636_ (.A(_0212_),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _1637_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .Y(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _1638_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1639_ (.A(_0214_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _1640_ (.A(_0212_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_1 _1641_ (.A(_0215_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _1642_ (.A(_0212_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _1643_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .Y(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _1644_ (.A(_0212_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _1645_ (.A(_0216_),
    .X(_0415_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(_0212_),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .Y(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _1648_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _1649_ (.A(_0217_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1650_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _1651_ (.A(_0218_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _1652_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_1 _1653_ (.A(_0219_),
    .X(_0414_));
 sky130_fd_sc_hd__inv_2 _1654_ (.A(_0212_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .Y(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _1656_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1657_ (.A(_0220_),
    .X(_0413_));
 sky130_fd_sc_hd__inv_2 _1658_ (.A(_0212_),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _1659_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .Y(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _1660_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _1661_ (.A(_0221_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _1662_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1663_ (.A(_0222_),
    .X(_0412_));
 sky130_fd_sc_hd__inv_2 _1664_ (.A(_0212_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .Y(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _1666_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_1 _1667_ (.A(_0223_),
    .X(_0411_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(_0212_),
    .Y(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _1669_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _1670_ (.A(_0224_),
    .X(_0799_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(_0165_),
    .Y(_0806_));
 sky130_fd_sc_hd__clkbuf_1 _1672_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .X(_0225_));
 sky130_fd_sc_hd__buf_1 _1673_ (.A(_0225_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _1674_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _1675_ (.A(_0226_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _1676_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _1677_ (.A(_0227_),
    .X(_0449_));
 sky130_fd_sc_hd__inv_2 _1678_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .Y(_0435_));
 sky130_fd_sc_hd__buf_6 _1679_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _1681_ (.A(_0229_),
    .X(_0445_));
 sky130_fd_sc_hd__inv_2 _1682_ (.A(_0228_),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _1683_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .Y(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(_0230_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _1686_ (.A(_0228_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(_0231_),
    .X(_0444_));
 sky130_fd_sc_hd__inv_2 _1688_ (.A(_0228_),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _1689_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .Y(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _1690_ (.A(_0228_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _1691_ (.A(_0232_),
    .X(_0443_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(_0228_),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .Y(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _1694_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _1695_ (.A(_0233_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _1696_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _1697_ (.A(_0234_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _1698_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_1 _1699_ (.A(_0235_),
    .X(_0442_));
 sky130_fd_sc_hd__inv_2 _1700_ (.A(_0228_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _1701_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .Y(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _1702_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(_0236_));
 sky130_fd_sc_hd__clkbuf_1 _1703_ (.A(_0236_),
    .X(_0441_));
 sky130_fd_sc_hd__inv_2 _1704_ (.A(_0228_),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_2 _1705_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .Y(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1706_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _1707_ (.A(_0237_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _1708_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _1709_ (.A(_0238_),
    .X(_0440_));
 sky130_fd_sc_hd__inv_2 _1710_ (.A(_0228_),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_2 _1711_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .Y(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _1712_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_1 _1713_ (.A(_0239_),
    .X(_0439_));
 sky130_fd_sc_hd__inv_2 _1714_ (.A(_0228_),
    .Y(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _1715_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _1716_ (.A(_0240_),
    .X(_0791_));
 sky130_fd_sc_hd__clkbuf_1 _1717_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .X(_0241_));
 sky130_fd_sc_hd__buf_1 _1718_ (.A(_0241_),
    .X(_0790_));
 sky130_fd_sc_hd__inv_2 _1719_ (.A(_0162_),
    .Y(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1720_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .X(_0242_));
 sky130_fd_sc_hd__buf_1 _1721_ (.A(_0242_),
    .X(_0824_));
 sky130_fd_sc_hd__inv_2 _1722_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .Y(_0549_));
 sky130_fd_sc_hd__clkbuf_1 _1723_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _1724_ (.A(_0243_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _1725_ (.A(_0162_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _1726_ (.A(_0244_),
    .X(_0556_));
 sky130_fd_sc_hd__inv_2 _1727_ (.A(_0162_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _1728_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .Y(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _1729_ (.A(_0162_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _1730_ (.A(_0245_),
    .X(_0555_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(_0162_),
    .Y(_0541_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .Y(_0550_));
 sky130_fd_sc_hd__clkbuf_1 _1733_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _1734_ (.A(_0246_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _1735_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _1736_ (.A(_0247_),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_1 _1737_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _1738_ (.A(_0248_),
    .X(_0554_));
 sky130_fd_sc_hd__inv_2 _1739_ (.A(_0162_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _1740_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .Y(_0545_));
 sky130_fd_sc_hd__clkbuf_1 _1741_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_1 _1742_ (.A(_0249_),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _1743_ (.A(_0162_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_2 _1744_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .Y(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _1745_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _1746_ (.A(_0250_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_1 _1748_ (.A(_0251_),
    .X(_0552_));
 sky130_fd_sc_hd__inv_2 _1749_ (.A(_0162_),
    .Y(_0538_));
 sky130_fd_sc_hd__inv_2 _1750_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .Y(_0544_));
 sky130_fd_sc_hd__clkbuf_1 _1751_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _1752_ (.A(_0252_),
    .X(_0551_));
 sky130_fd_sc_hd__inv_2 _1753_ (.A(_0162_),
    .Y(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1754_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _1755_ (.A(_0253_),
    .X(_0825_));
 sky130_fd_sc_hd__inv_2 _1756_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _1757_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .Y(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _1758_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _1759_ (.A(_0254_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _1760_ (.A(_0096_),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_1 _1761_ (.A(_0255_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _1762_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .X(_0256_));
 sky130_fd_sc_hd__buf_1 _1763_ (.A(_0256_),
    .X(_0858_));
 sky130_fd_sc_hd__inv_2 _1764_ (.A(_0096_),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .Y(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _1766_ (.A(_0096_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_1 _1767_ (.A(_0257_),
    .X(_0667_));
 sky130_fd_sc_hd__inv_2 _1768_ (.A(_0096_),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _1769_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .Y(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _1770_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .X(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _1771_ (.A(_0258_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _1772_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _1773_ (.A(_0259_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _1774_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _1775_ (.A(_0260_),
    .X(_0666_));
 sky130_fd_sc_hd__inv_2 _1776_ (.A(_0096_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _1777_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .Y(_0657_));
 sky130_fd_sc_hd__clkbuf_1 _1778_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_1 _1779_ (.A(_0261_),
    .X(_0665_));
 sky130_fd_sc_hd__inv_2 _1780_ (.A(_0096_),
    .Y(_0651_));
 sky130_fd_sc_hd__inv_2 _1781_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .Y(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _1782_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _1783_ (.A(_0262_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _1784_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_1 _1785_ (.A(_0263_),
    .X(_0664_));
 sky130_fd_sc_hd__inv_2 _1786_ (.A(_0096_),
    .Y(_0650_));
 sky130_fd_sc_hd__inv_2 _1787_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .Y(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1788_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(_0264_),
    .X(_0663_));
 sky130_fd_sc_hd__inv_2 _1790_ (.A(_0096_),
    .Y(_0649_));
 sky130_fd_sc_hd__clkbuf_1 _1791_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _1792_ (.A(_0265_),
    .X(_0859_));
 sky130_fd_sc_hd__inv_2 _1793_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .Y(_0855_));
 sky130_fd_sc_hd__inv_2 _1794_ (.A(_0028_),
    .Y(_0766_));
 sky130_fd_sc_hd__clkbuf_1 _1795_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .X(_0266_));
 sky130_fd_sc_hd__buf_1 _1796_ (.A(_0266_),
    .X(_0892_));
 sky130_fd_sc_hd__inv_2 _1797_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .Y(_0770_));
 sky130_fd_sc_hd__clkbuf_1 _1798_ (.A(_0028_),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_1 _1799_ (.A(_0267_),
    .X(_0779_));
 sky130_fd_sc_hd__inv_2 _1800_ (.A(_0028_),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_2 _1801_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .Y(_0774_));
 sky130_fd_sc_hd__clkbuf_1 _1802_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _1803_ (.A(_0268_),
    .X(_0786_));
 sky130_fd_sc_hd__clkbuf_1 _1804_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_1 _1805_ (.A(_0269_),
    .X(_0783_));
 sky130_fd_sc_hd__clkbuf_1 _1806_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _1807_ (.A(_0270_),
    .X(_0778_));
 sky130_fd_sc_hd__inv_2 _1808_ (.A(_0028_),
    .Y(_0764_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .Y(_0769_));
 sky130_fd_sc_hd__clkbuf_1 _1810_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _1811_ (.A(_0271_),
    .X(_0777_));
 sky130_fd_sc_hd__inv_2 _1812_ (.A(_0028_),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_2 _1813_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .Y(_0772_));
 sky130_fd_sc_hd__clkbuf_1 _1814_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_1 _1815_ (.A(_0272_),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_1 _1816_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _1817_ (.A(_0273_),
    .X(_0776_));
 sky130_fd_sc_hd__inv_2 _1818_ (.A(_0028_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _1819_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .Y(_0768_));
 sky130_fd_sc_hd__clkbuf_1 _1820_ (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _1821_ (.A(_0274_),
    .X(_0775_));
 sky130_fd_sc_hd__inv_2 _1822_ (.A(_0028_),
    .Y(_0761_));
 sky130_fd_sc_hd__clkbuf_1 _1823_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _1824_ (.A(_0275_),
    .X(_0893_));
 sky130_fd_sc_hd__inv_2 _1825_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .Y(_0889_));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(_0176_),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(_0176_),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _1828_ (.A(_0176_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _1829_ (.A(_0176_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(_0176_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _1831_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__inv_2 _1832_ (.A(net12),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(net8),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _1834_ (.A(net1),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _1835_ (.A(net5),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _1836_ (.A(net13),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _1837_ (.A(net9),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _1838_ (.A(net2),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(net6),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(net14),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _1841_ (.A(net10),
    .Y(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _1842_ (.A(net27),
    .Y(net18));
 sky130_fd_sc_hd__inv_2 _1843_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _1844_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _1845_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _1846_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _1848_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _1849_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _1853_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _1854_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _1855_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ));
 sky130_fd_sc_hd__inv_2 _1857_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ));
 sky130_fd_sc_hd__inv_2 _1858_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__inv_2 _1860_ (.A(net23),
    .Y(net19));
 sky130_fd_sc_hd__inv_2 _1861_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _1863_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _1864_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _1865_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _1866_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _1867_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _1869_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _1870_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _1871_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ));
 sky130_fd_sc_hd__inv_2 _1874_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ));
 sky130_fd_sc_hd__inv_2 _1875_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ));
 sky130_fd_sc_hd__inv_2 _1876_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ));
 sky130_fd_sc_hd__inv_2 _1877_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__inv_2 _1878_ (.A(net20),
    .Y(net17));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _1880_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _1881_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _1882_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _1883_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _1884_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _1885_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _1886_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _1888_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _1889_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _1890_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _1891_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ));
 sky130_fd_sc_hd__inv_2 _1892_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ));
 sky130_fd_sc_hd__inv_2 _1893_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ));
 sky130_fd_sc_hd__inv_2 _1894_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ));
 sky130_fd_sc_hd__inv_2 _1895_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ));
 sky130_fd_sc_hd__inv_2 _1896_ (.A(net24),
    .Y(net15));
 sky130_fd_sc_hd__inv_2 _1897_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _1898_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _1899_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _1900_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _1901_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _1902_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _1903_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _1904_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _1905_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _1906_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ));
 sky130_fd_sc_hd__inv_2 _1907_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ));
 sky130_fd_sc_hd__inv_2 _1908_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ));
 sky130_fd_sc_hd__inv_2 _1909_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ));
 sky130_fd_sc_hd__inv_2 _1910_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ));
 sky130_fd_sc_hd__inv_2 _1911_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ));
 sky130_fd_sc_hd__inv_2 _1912_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .Y(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ));
 sky130_fd_sc_hd__inv_2 _1913_ (.A(_0176_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _1914_ (.A(net4),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1915_ (.A(net4),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1916_ (.A(net4),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1917_ (.A(net4),
    .Y(_0011_));
 sky130_fd_sc_hd__dfxtp_1 _1918_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net68),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _1919_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net136),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1920_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net99),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1921_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net100),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net116),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net107),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1924_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net119),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1925_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net111),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net98),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1927_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net127),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net69),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net85),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net91),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net106),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net151),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net3),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net205),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _1935_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net79),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfbbn_1 _1936_ (.CLK_N(_0002_),
    .D(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(_0000_),
    .SET_B(_0001_),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfxtp_1 _1937_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net146),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1938_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net176),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net194),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net175),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net139),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1942_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net152),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net182),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net174),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1945_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net149),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1946_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net183),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net192),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net170),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net203),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1950_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net156),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net200),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1952_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net186),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net76),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1954_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net165),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net207),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net177),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net140),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1958_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net187),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net197),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1960_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net190),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1961_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net148),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1962_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net166),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1963_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net196),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1964_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net159),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1965_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net206),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1966_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net169),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1967_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net201),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1968_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net178),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1969_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net74),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1970_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net162),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1971_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net191),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1972_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net180),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1973_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net147),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1974_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net179),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1975_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net202),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1976_ (.CLK(clknet_4_3_0_prog_clk),
    .D(net171),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1977_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net155),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1978_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net173),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1979_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net198),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1980_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net158),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1981_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net154),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1982_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net163),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1983_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net185),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1984_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net181),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1985_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net77),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1986_ (.CLK(clknet_4_9_0_prog_clk),
    .D(net160),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1987_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net164),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1988_ (.CLK(clknet_4_10_0_prog_clk),
    .D(net189),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1989_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net129),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1990_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net168),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1991_ (.CLK(clknet_4_12_0_prog_clk),
    .D(net195),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1992_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net161),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1993_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net150),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1994_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net167),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1995_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net188),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1996_ (.CLK(clknet_4_11_0_prog_clk),
    .D(net184),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1997_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net94),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _1998_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net153),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _1999_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net193),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2000_ (.CLK(clknet_4_14_0_prog_clk),
    .D(net172),
    .Q(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2001_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net89),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _2002_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net87),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2003_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net125),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2004_ (.CLK(clknet_4_15_0_prog_clk),
    .D(net72),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2005_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net78),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2006_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net80),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2007_ (.CLK(clknet_4_13_0_prog_clk),
    .D(net92),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2008_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net104),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2009_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net109),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2010_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net132),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2011_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net130),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2012_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net126),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2013_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net128),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2014_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net101),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2015_ (.CLK(clknet_4_7_0_prog_clk),
    .D(net70),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2016_ (.CLK(clknet_4_6_0_prog_clk),
    .D(net133),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfbbn_1 _2017_ (.CLK_N(_0005_),
    .D(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(_0003_),
    .SET_B(_0004_),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfxtp_1 _2018_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net84),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2019_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net138),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _2020_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net93),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _2021_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net88),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2022_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net123),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2023_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net97),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2024_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net102),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2025_ (.CLK(clknet_4_5_0_prog_clk),
    .D(net71),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2026_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net81),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2027_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net108),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2028_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net86),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2029_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net95),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2030_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net83),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2031_ (.CLK(clknet_4_4_0_prog_clk),
    .D(net82),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2032_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net113),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2033_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net112),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2034_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net110),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2035_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net157),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfbbn_1 _2036_ (.CLK_N(_0008_),
    .D(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(_0006_),
    .SET_B(_0007_),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfxtp_1 _2037_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net90),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2038_ (.CLK(clknet_4_1_0_prog_clk),
    .D(net137),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _2039_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net96),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 _2040_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net103),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2041_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net114),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2042_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net122),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2043_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net121),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2044_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net115),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2045_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net117),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2046_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net135),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2047_ (.CLK(clknet_4_0_0_prog_clk),
    .D(net73),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2048_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net120),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2049_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net124),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2050_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net118),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2051_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net131),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2052_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net105),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2053_ (.CLK(clknet_4_2_0_prog_clk),
    .D(net75),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ));
 sky130_fd_sc_hd__dfxtp_1 _2054_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net141),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ));
 sky130_fd_sc_hd__dfbbn_1 _2055_ (.CLK_N(_0011_),
    .D(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.direct_interc_4_.in ),
    .RESET_B(_0009_),
    .SET_B(_0010_),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.Q ),
    .Q_N(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfxtp_1 _2056_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net134),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2057_ (.CLK(clknet_4_8_0_prog_clk),
    .D(net204),
    .Q(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ));
 sky130_fd_sc_hd__ebufn_1 _2078_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ),
    .TE_B(_0324_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2079_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ),
    .TE_B(_0325_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2080_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ),
    .TE_B(_0326_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2081_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ),
    .TE_B(_0327_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2082_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ),
    .TE_B(_0328_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2083_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ),
    .TE_B(_0329_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2084_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ),
    .TE_B(_0330_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2085_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ),
    .TE_B(_0331_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2086_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ),
    .TE_B(_0332_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2087_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ),
    .TE_B(_0333_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2088_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ),
    .TE_B(_0334_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2089_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ),
    .TE_B(_0335_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2090_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ),
    .TE_B(_0336_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2091_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ),
    .TE_B(_0337_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2092_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ),
    .TE_B(_0338_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_8 _2093_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0339_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2094_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0340_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2095_ (.A(net47),
    .TE_B(_0341_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2096_ (.A(net42),
    .TE_B(_0342_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2097_ (.A(net39),
    .TE_B(_0343_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2098_ (.A(net35),
    .TE_B(_0344_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2099_ (.A(net30),
    .TE_B(_0345_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2100_ (.A(net24),
    .TE_B(_0346_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2101_ (.A(net23),
    .TE_B(_0347_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2102_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0348_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2103_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0349_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2104_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0350_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2105_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0351_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2106_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0352_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2107_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0353_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2108_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0354_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2109_ (.A(net45),
    .TE_B(_0355_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2110_ (.A(net40),
    .TE_B(_0356_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2111_ (.A(net37),
    .TE_B(_0357_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2112_ (.A(net33),
    .TE_B(_0358_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2113_ (.A(net29),
    .TE_B(_0359_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2114_ (.A(net20),
    .TE_B(_0360_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2115_ (.A(net26),
    .TE_B(_0361_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2116_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0362_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2117_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0363_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2118_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0364_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2119_ (.A(net48),
    .TE_B(_0365_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2119__48 (.HI(net48));
 sky130_fd_sc_hd__ebufn_1 _2120_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0366_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2121_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0367_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2122_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0368_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2123_ (.A(net47),
    .TE_B(_0369_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2124_ (.A(net42),
    .TE_B(_0370_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2125_ (.A(net39),
    .TE_B(_0371_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2126_ (.A(net35),
    .TE_B(_0372_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2127_ (.A(net31),
    .TE_B(_0373_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2128_ (.A(net24),
    .TE_B(_0374_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2129_ (.A(net23),
    .TE_B(_0375_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2130_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0376_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2131_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0377_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2132_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0378_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2133_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0379_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2134_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0380_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2135_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0381_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2136_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0382_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2137_ (.A(net45),
    .TE_B(_0383_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2138_ (.A(net40),
    .TE_B(_0384_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2139_ (.A(net37),
    .TE_B(_0385_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2140_ (.A(net33),
    .TE_B(_0386_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2141_ (.A(net29),
    .TE_B(_0387_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2142_ (.A(net20),
    .TE_B(_0388_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2143_ (.A(net27),
    .TE_B(_0389_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2144_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0390_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2145_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0391_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2146_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0392_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2147_ (.A(net49),
    .TE_B(_0393_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2147__49 (.HI(net49));
 sky130_fd_sc_hd__ebufn_1 _2148_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0394_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2149_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0395_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2150_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0396_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2151_ (.A(net47),
    .TE_B(_0397_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2152_ (.A(net42),
    .TE_B(_0398_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2153_ (.A(net38),
    .TE_B(_0399_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2154_ (.A(net34),
    .TE_B(_0400_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2155_ (.A(net30),
    .TE_B(_0401_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2156_ (.A(net25),
    .TE_B(_0402_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2157_ (.A(net23),
    .TE_B(_0403_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2158_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0404_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2159_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0405_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2160_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0406_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2161_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0407_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2162_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0408_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2163_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0409_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2164_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0410_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2165_ (.A(net45),
    .TE_B(_0411_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2166_ (.A(net40),
    .TE_B(_0412_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2167_ (.A(net36),
    .TE_B(_0413_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2168_ (.A(net32),
    .TE_B(_0414_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2169_ (.A(net28),
    .TE_B(_0415_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2170_ (.A(net21),
    .TE_B(_0416_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2171_ (.A(net26),
    .TE_B(_0417_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2172_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0418_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2173_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0419_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2174_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0420_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2175_ (.A(net50),
    .TE_B(_0421_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2175__50 (.HI(net50));
 sky130_fd_sc_hd__ebufn_2 _2176_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0422_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2177_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0423_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2178_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0424_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_2 _2179_ (.A(net46),
    .TE_B(_0425_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2180_ (.A(net42),
    .TE_B(_0426_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2181_ (.A(net38),
    .TE_B(_0427_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2182_ (.A(net34),
    .TE_B(_0428_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2183_ (.A(net30),
    .TE_B(_0429_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2184_ (.A(net25),
    .TE_B(_0430_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2185_ (.A(net22),
    .TE_B(_0431_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2186_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0432_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2187_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0433_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2188_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0434_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2189_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0435_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2190_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0436_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2191_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0437_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2192_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0438_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2193_ (.A(net44),
    .TE_B(_0439_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2194_ (.A(net40),
    .TE_B(_0440_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2195_ (.A(net36),
    .TE_B(_0441_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2196_ (.A(net32),
    .TE_B(_0442_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2197_ (.A(net28),
    .TE_B(_0443_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2198_ (.A(net20),
    .TE_B(_0444_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2199_ (.A(net26),
    .TE_B(_0445_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2200_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0446_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2201_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0447_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2202_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0448_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2203_ (.A(net51),
    .TE_B(_0449_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2203__51 (.HI(net51));
 sky130_fd_sc_hd__ebufn_4 _2204_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0450_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2205_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0451_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2206_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0452_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2207_ (.A(net46),
    .TE_B(_0453_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2208_ (.A(net42),
    .TE_B(_0454_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2209_ (.A(net38),
    .TE_B(_0455_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2210_ (.A(net34),
    .TE_B(_0456_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2211_ (.A(net30),
    .TE_B(_0457_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2212_ (.A(net25),
    .TE_B(_0458_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2213_ (.A(net22),
    .TE_B(_0459_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2214_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0460_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2215_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0461_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2216_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0462_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2217_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0463_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2218_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0464_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2219_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0465_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2220_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0466_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2221_ (.A(net44),
    .TE_B(_0467_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2222_ (.A(net40),
    .TE_B(_0468_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2223_ (.A(net36),
    .TE_B(_0469_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2224_ (.A(net32),
    .TE_B(_0470_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2225_ (.A(net28),
    .TE_B(_0471_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2226_ (.A(net20),
    .TE_B(_0472_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2227_ (.A(net26),
    .TE_B(_0473_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2228_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0474_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2229_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0475_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2230_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0476_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2231_ (.A(net52),
    .TE_B(_0477_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2231__52 (.HI(net52));
 sky130_fd_sc_hd__ebufn_1 _2232_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0478_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2233_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0479_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2234_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0480_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2235_ (.A(net46),
    .TE_B(_0481_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2236_ (.A(net42),
    .TE_B(_0482_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2237_ (.A(net38),
    .TE_B(_0483_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2238_ (.A(net34),
    .TE_B(_0484_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2239_ (.A(net30),
    .TE_B(_0485_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2240_ (.A(net25),
    .TE_B(_0486_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2241_ (.A(net22),
    .TE_B(_0487_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2242_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0488_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2243_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0489_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2244_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0490_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2245_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0491_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2246_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0492_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2247_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0493_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2248_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0494_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2249_ (.A(net44),
    .TE_B(_0495_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2250_ (.A(net40),
    .TE_B(_0496_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2251_ (.A(net36),
    .TE_B(_0497_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2252_ (.A(net32),
    .TE_B(_0498_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2253_ (.A(net28),
    .TE_B(_0499_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2254_ (.A(net20),
    .TE_B(_0500_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2255_ (.A(net26),
    .TE_B(_0501_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2256_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0502_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2257_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0503_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2258_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0504_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2259_ (.A(net53),
    .TE_B(_0505_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2259__53 (.HI(net53));
 sky130_fd_sc_hd__ebufn_1 _2260_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0506_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2261_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0507_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2262_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0508_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2263_ (.A(net46),
    .TE_B(_0509_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2264_ (.A(net42),
    .TE_B(_0510_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2265_ (.A(net38),
    .TE_B(_0511_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2266_ (.A(net34),
    .TE_B(_0512_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2267_ (.A(net30),
    .TE_B(_0513_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2268_ (.A(net24),
    .TE_B(_0514_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2269_ (.A(net23),
    .TE_B(_0515_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2270_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0516_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2271_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0517_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2272_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0518_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2273_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0519_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2274_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0520_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2275_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0521_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2276_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0522_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2277_ (.A(net44),
    .TE_B(_0523_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2278_ (.A(net40),
    .TE_B(_0524_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2279_ (.A(net36),
    .TE_B(_0525_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2280_ (.A(net32),
    .TE_B(_0526_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2281_ (.A(net28),
    .TE_B(_0527_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2282_ (.A(net20),
    .TE_B(_0528_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2283_ (.A(net26),
    .TE_B(_0529_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2284_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0530_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2285_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0531_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2286_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0532_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2287_ (.A(net54),
    .TE_B(_0533_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2287__54 (.HI(net54));
 sky130_fd_sc_hd__ebufn_1 _2288_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0534_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2289_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0535_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2290_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0536_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2291_ (.A(net46),
    .TE_B(_0537_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2292_ (.A(net42),
    .TE_B(_0538_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2293_ (.A(net38),
    .TE_B(_0539_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2294_ (.A(net34),
    .TE_B(_0540_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2295_ (.A(net30),
    .TE_B(_0541_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2296_ (.A(net24),
    .TE_B(_0542_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2297_ (.A(net22),
    .TE_B(_0543_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2298_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0544_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2299_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0545_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2300_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0546_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2301_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0547_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2302_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0548_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2303_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0549_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2304_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0550_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2305_ (.A(net44),
    .TE_B(_0551_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2306_ (.A(net40),
    .TE_B(_0552_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2307_ (.A(net36),
    .TE_B(_0553_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2308_ (.A(net32),
    .TE_B(_0554_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2309_ (.A(net28),
    .TE_B(_0555_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2310_ (.A(net20),
    .TE_B(_0556_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2311_ (.A(net26),
    .TE_B(_0557_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2312_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0558_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2313_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0559_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2314_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0560_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2315_ (.A(net55),
    .TE_B(_0561_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2315__55 (.HI(net55));
 sky130_fd_sc_hd__ebufn_1 _2316_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0562_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2317_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0563_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2318_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0564_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2319_ (.A(net46),
    .TE_B(_0565_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2320_ (.A(net42),
    .TE_B(_0566_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2321_ (.A(net38),
    .TE_B(_0567_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2322_ (.A(net34),
    .TE_B(_0568_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2323_ (.A(net30),
    .TE_B(_0569_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2324_ (.A(net24),
    .TE_B(_0570_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2325_ (.A(net22),
    .TE_B(_0571_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2326_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0572_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2327_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0573_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2328_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0574_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2329_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0575_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2330_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0576_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2331_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0577_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2332_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0578_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2333_ (.A(net44),
    .TE_B(_0579_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2334_ (.A(net40),
    .TE_B(_0580_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2335_ (.A(net36),
    .TE_B(_0581_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2336_ (.A(net32),
    .TE_B(_0582_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2337_ (.A(net28),
    .TE_B(_0583_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2338_ (.A(net20),
    .TE_B(_0584_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2339_ (.A(net26),
    .TE_B(_0585_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2340_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0586_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2341_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0587_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2342_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0588_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2343_ (.A(net56),
    .TE_B(_0589_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2343__56 (.HI(net56));
 sky130_fd_sc_hd__ebufn_1 _2344_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0590_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2345_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0591_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2346_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0592_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2347_ (.A(net46),
    .TE_B(_0593_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2348_ (.A(net42),
    .TE_B(_0594_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2349_ (.A(net38),
    .TE_B(_0595_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2350_ (.A(net34),
    .TE_B(_0596_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2351_ (.A(net30),
    .TE_B(_0597_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2352_ (.A(net24),
    .TE_B(_0598_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2353_ (.A(net22),
    .TE_B(_0599_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2354_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0600_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2355_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0601_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2356_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0602_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2357_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0603_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2358_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0604_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2359_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0605_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2360_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0606_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2361_ (.A(net44),
    .TE_B(_0607_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2362_ (.A(net40),
    .TE_B(_0608_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2363_ (.A(net36),
    .TE_B(_0609_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2364_ (.A(net32),
    .TE_B(_0610_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2365_ (.A(net28),
    .TE_B(_0611_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2366_ (.A(net20),
    .TE_B(_0612_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2367_ (.A(net26),
    .TE_B(_0613_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2368_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0614_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2369_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0615_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2370_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0616_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2371_ (.A(net57),
    .TE_B(_0617_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2371__57 (.HI(net57));
 sky130_fd_sc_hd__ebufn_1 _2372_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0618_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2373_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0619_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2374_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0620_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2375_ (.A(net46),
    .TE_B(_0621_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2376_ (.A(net43),
    .TE_B(_0622_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2377_ (.A(net38),
    .TE_B(_0623_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2378_ (.A(net34),
    .TE_B(_0624_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2379_ (.A(net30),
    .TE_B(_0625_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2380_ (.A(net24),
    .TE_B(_0626_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2381_ (.A(net22),
    .TE_B(_0627_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2382_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0628_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2383_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0629_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2384_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0630_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2385_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0631_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2386_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0632_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2387_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0633_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2388_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0634_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2389_ (.A(net44),
    .TE_B(_0635_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2390_ (.A(net41),
    .TE_B(_0636_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2391_ (.A(net36),
    .TE_B(_0637_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2392_ (.A(net32),
    .TE_B(_0638_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2393_ (.A(net28),
    .TE_B(_0639_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2394_ (.A(net21),
    .TE_B(_0640_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2395_ (.A(net26),
    .TE_B(_0641_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2396_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0642_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2397_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0643_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2398_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0644_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2399_ (.A(net58),
    .TE_B(_0645_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2399__58 (.HI(net58));
 sky130_fd_sc_hd__ebufn_1 _2400_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0646_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2401_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0647_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2402_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0648_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2403_ (.A(net46),
    .TE_B(_0649_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2404_ (.A(net43),
    .TE_B(_0650_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2405_ (.A(net38),
    .TE_B(_0651_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2406_ (.A(net35),
    .TE_B(_0652_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2407_ (.A(net31),
    .TE_B(_0653_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2408_ (.A(net24),
    .TE_B(_0654_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2409_ (.A(net23),
    .TE_B(_0655_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2410_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0656_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2411_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0657_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2412_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0658_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2413_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0659_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2414_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0660_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2415_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0661_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2416_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0662_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2417_ (.A(net44),
    .TE_B(_0663_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2418_ (.A(net41),
    .TE_B(_0664_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2419_ (.A(net37),
    .TE_B(_0665_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2420_ (.A(net33),
    .TE_B(_0666_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2421_ (.A(net29),
    .TE_B(_0667_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2422_ (.A(net21),
    .TE_B(_0668_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2423_ (.A(net27),
    .TE_B(_0669_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2424_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0670_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2425_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0671_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2426_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0672_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2427_ (.A(net59),
    .TE_B(_0673_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2427__59 (.HI(net59));
 sky130_fd_sc_hd__ebufn_2 _2428_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0674_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2429_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0675_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2430_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0676_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2431_ (.A(net46),
    .TE_B(_0677_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2432_ (.A(net43),
    .TE_B(_0678_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2433_ (.A(net39),
    .TE_B(_0679_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2434_ (.A(net35),
    .TE_B(_0680_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2435_ (.A(net31),
    .TE_B(_0681_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2436_ (.A(net24),
    .TE_B(_0682_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2437_ (.A(net22),
    .TE_B(_0683_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2438_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0684_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2439_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0685_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2440_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0686_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2441_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0687_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2442_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0688_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2443_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0689_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2444_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0690_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2445_ (.A(net44),
    .TE_B(_0691_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2446_ (.A(net41),
    .TE_B(_0692_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2447_ (.A(net37),
    .TE_B(_0693_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2448_ (.A(net33),
    .TE_B(_0694_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2449_ (.A(net29),
    .TE_B(_0695_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2450_ (.A(net21),
    .TE_B(_0696_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2451_ (.A(net27),
    .TE_B(_0697_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2452_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0698_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2453_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0699_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _2454_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0700_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2455_ (.A(net60),
    .TE_B(_0701_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2455__60 (.HI(net60));
 sky130_fd_sc_hd__ebufn_1 _2456_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0702_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2457_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0703_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2458_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0704_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.out ));
 sky130_fd_sc_hd__ebufn_1 _2459_ (.A(net47),
    .TE_B(_0705_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2460_ (.A(net43),
    .TE_B(_0706_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2461_ (.A(net39),
    .TE_B(_0707_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2462_ (.A(net34),
    .TE_B(_0708_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2463_ (.A(net31),
    .TE_B(_0709_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2464_ (.A(net25),
    .TE_B(_0710_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2465_ (.A(net22),
    .TE_B(_0711_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2466_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0712_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2467_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0713_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2468_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0714_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2469_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0715_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2470_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0716_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2471_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0717_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2472_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0718_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2473_ (.A(net45),
    .TE_B(_0719_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2474_ (.A(net41),
    .TE_B(_0720_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2475_ (.A(net37),
    .TE_B(_0721_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2476_ (.A(net33),
    .TE_B(_0722_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2477_ (.A(net28),
    .TE_B(_0723_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2478_ (.A(net21),
    .TE_B(_0724_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2479_ (.A(net27),
    .TE_B(_0725_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2480_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0726_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2481_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0727_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2482_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0728_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2483_ (.A(net61),
    .TE_B(_0729_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2483__61 (.HI(net61));
 sky130_fd_sc_hd__ebufn_1 _2484_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0730_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2485_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0731_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2486_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0732_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.out ));
 sky130_fd_sc_hd__ebufn_1 _2487_ (.A(net47),
    .TE_B(_0733_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2488_ (.A(net43),
    .TE_B(_0734_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2489_ (.A(net39),
    .TE_B(_0735_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2490_ (.A(net35),
    .TE_B(_0736_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2491_ (.A(net31),
    .TE_B(_0737_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2492_ (.A(net25),
    .TE_B(_0738_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2493_ (.A(net22),
    .TE_B(_0739_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2494_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0740_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2495_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0741_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2496_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0742_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2497_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0743_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2498_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0744_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2499_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0745_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2500_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0746_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2501_ (.A(net45),
    .TE_B(_0747_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2502_ (.A(net41),
    .TE_B(_0748_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2503_ (.A(net36),
    .TE_B(_0749_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2504_ (.A(net32),
    .TE_B(_0750_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2505_ (.A(net29),
    .TE_B(_0751_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2506_ (.A(net21),
    .TE_B(_0752_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2507_ (.A(net27),
    .TE_B(_0753_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2508_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0754_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2509_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0755_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2510_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0756_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2511_ (.A(net62),
    .TE_B(_0757_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2511__62 (.HI(net62));
 sky130_fd_sc_hd__ebufn_1 _2512_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0758_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2513_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0759_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2514_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0760_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.out ));
 sky130_fd_sc_hd__ebufn_1 _2515_ (.A(net47),
    .TE_B(_0761_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2516_ (.A(net43),
    .TE_B(_0762_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2517_ (.A(net39),
    .TE_B(_0763_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2518_ (.A(net35),
    .TE_B(_0764_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2519_ (.A(net31),
    .TE_B(_0765_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2520_ (.A(net25),
    .TE_B(_0766_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2521_ (.A(net23),
    .TE_B(_0767_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2522_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0768_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2523_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .TE_B(_0769_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2524_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out ),
    .TE_B(_0770_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2525_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out ),
    .TE_B(_0771_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2526_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_0772_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2527_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_0773_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2528_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_0774_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2529_ (.A(net45),
    .TE_B(_0775_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2530_ (.A(net41),
    .TE_B(_0776_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2531_ (.A(net37),
    .TE_B(_0777_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2532_ (.A(net33),
    .TE_B(_0778_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2533_ (.A(net29),
    .TE_B(_0779_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2534_ (.A(net21),
    .TE_B(_0780_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2535_ (.A(net27),
    .TE_B(_0781_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2536_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_0782_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2537_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .TE_B(_0783_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2538_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.out ),
    .TE_B(_0784_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2539_ (.A(net63),
    .TE_B(_0785_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2539__63 (.HI(net63));
 sky130_fd_sc_hd__ebufn_1 _2540_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_0786_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _2541_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_0787_),
    .Z(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2542_ (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_0788_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2543_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0789_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2544_ (.A(net64),
    .TE_B(_0790_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2544__64 (.HI(net64));
 sky130_fd_sc_hd__ebufn_1 _2545_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ),
    .TE_B(_0791_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2546_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ),
    .TE_B(_0792_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2547_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ),
    .TE_B(_0793_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2548_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ),
    .TE_B(_0794_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2549_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ),
    .TE_B(_0795_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2550_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ),
    .TE_B(_0796_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2551_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ),
    .TE_B(_0797_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2552_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ),
    .TE_B(_0798_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2553_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ),
    .TE_B(_0799_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2554_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ),
    .TE_B(_0800_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2555_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ),
    .TE_B(_0801_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2556_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ),
    .TE_B(_0802_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2557_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ),
    .TE_B(_0803_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2558_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ),
    .TE_B(_0804_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2559_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ),
    .TE_B(_0805_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2560_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ),
    .TE_B(_0806_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2561_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ),
    .TE_B(_0807_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2562_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ),
    .TE_B(_0808_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2563_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ),
    .TE_B(_0809_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2564_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ),
    .TE_B(_0810_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2565_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ),
    .TE_B(_0811_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2566_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ),
    .TE_B(_0812_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2567_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ),
    .TE_B(_0813_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2568_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ),
    .TE_B(_0814_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2569_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ),
    .TE_B(_0815_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2570_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ),
    .TE_B(_0816_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_2 _2571_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ),
    .TE_B(_0817_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2572_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ),
    .TE_B(_0818_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_4 _2573_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ),
    .TE_B(_0819_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_8 _2574_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ),
    .TE_B(_0820_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2575_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0821_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2576_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0822_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2577_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0823_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2578_ (.A(net65),
    .TE_B(_0824_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2578__65 (.HI(net65));
 sky130_fd_sc_hd__ebufn_1 _2579_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ),
    .TE_B(_0825_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2580_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ),
    .TE_B(_0826_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2581_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ),
    .TE_B(_0827_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2582_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ),
    .TE_B(_0828_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2583_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ),
    .TE_B(_0829_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2584_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ),
    .TE_B(_0830_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2585_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ),
    .TE_B(_0831_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2586_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ),
    .TE_B(_0832_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2587_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ),
    .TE_B(_0833_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2588_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ),
    .TE_B(_0834_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2589_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ),
    .TE_B(_0835_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2590_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ),
    .TE_B(_0836_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2591_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ),
    .TE_B(_0837_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2592_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ),
    .TE_B(_0838_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2593_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ),
    .TE_B(_0839_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2594_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ),
    .TE_B(_0840_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2595_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ),
    .TE_B(_0841_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2596_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ),
    .TE_B(_0842_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2597_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ),
    .TE_B(_0843_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2598_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ),
    .TE_B(_0844_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2599_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ),
    .TE_B(_0845_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2600_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ),
    .TE_B(_0846_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2601_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ),
    .TE_B(_0847_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2602_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ),
    .TE_B(_0848_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2603_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ),
    .TE_B(_0849_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2604_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ),
    .TE_B(_0850_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2605_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ),
    .TE_B(_0851_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2606_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ),
    .TE_B(_0852_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2607_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ),
    .TE_B(_0853_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2608_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ),
    .TE_B(_0854_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2609_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0855_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2610_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0856_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2611_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0857_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2612_ (.A(net66),
    .TE_B(_0858_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2612__66 (.HI(net66));
 sky130_fd_sc_hd__ebufn_1 _2613_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ),
    .TE_B(_0859_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2614_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ),
    .TE_B(_0860_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2615_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ),
    .TE_B(_0861_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2616_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ),
    .TE_B(_0862_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2617_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ),
    .TE_B(_0863_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2618_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ),
    .TE_B(_0864_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2619_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ),
    .TE_B(_0865_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2620_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ),
    .TE_B(_0866_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2621_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ),
    .TE_B(_0867_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2622_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ),
    .TE_B(_0868_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2623_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ),
    .TE_B(_0869_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2624_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ),
    .TE_B(_0870_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2625_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ),
    .TE_B(_0871_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2626_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ),
    .TE_B(_0872_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2627_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ),
    .TE_B(_0873_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2628_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.out ),
    .TE_B(_0874_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2629_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.out ),
    .TE_B(_0875_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2630_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.out ),
    .TE_B(_0876_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2631_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.out ),
    .TE_B(_0877_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2632_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.out ),
    .TE_B(_0878_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2633_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.out ),
    .TE_B(_0879_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2634_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.out ),
    .TE_B(_0880_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2635_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.out ),
    .TE_B(_0881_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2636_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ),
    .TE_B(_0882_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2637_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ),
    .TE_B(_0883_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2638_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ),
    .TE_B(_0884_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2639_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ),
    .TE_B(_0885_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2640_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ),
    .TE_B(_0886_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2641_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ),
    .TE_B(_0887_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2642_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ),
    .TE_B(_0888_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__ebufn_1 _2643_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0889_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_8 _2644_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_0890_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2645_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0891_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_4 _2646_ (.A(net67),
    .TE_B(_0892_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _2646__67 (.HI(net67));
 sky130_fd_sc_hd__ebufn_1 _2647_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.out ),
    .TE_B(_0893_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _2648_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.out ),
    .TE_B(_0894_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _2649_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.out ),
    .TE_B(_0895_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _2650_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.out ),
    .TE_B(_0896_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_3_out ));
 sky130_fd_sc_hd__ebufn_1 _2651_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.out ),
    .TE_B(_0897_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ));
 sky130_fd_sc_hd__ebufn_1 _2652_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.out ),
    .TE_B(_0898_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_5_out ));
 sky130_fd_sc_hd__ebufn_1 _2653_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.out ),
    .TE_B(_0899_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ));
 sky130_fd_sc_hd__ebufn_1 _2654_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.out ),
    .TE_B(_0900_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_7_out ));
 sky130_fd_sc_hd__ebufn_1 _2655_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_0_out ),
    .TE_B(_0901_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ));
 sky130_fd_sc_hd__ebufn_1 _2656_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_2_out ),
    .TE_B(_0902_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_9_out ));
 sky130_fd_sc_hd__ebufn_1 _2657_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_4_out ),
    .TE_B(_0903_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ));
 sky130_fd_sc_hd__ebufn_1 _2658_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_6_out ),
    .TE_B(_0904_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_11_out ));
 sky130_fd_sc_hd__ebufn_1 _2659_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_8_out ),
    .TE_B(_0905_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ));
 sky130_fd_sc_hd__ebufn_1 _2660_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_10_out ),
    .TE_B(_0906_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_13_out ));
 sky130_fd_sc_hd__ebufn_2 _2661_ (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.lut4_mux_basis_input2_mem1_12_out ),
    .TE_B(_0907_),
    .Z(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_0_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_10_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_11_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_12_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_13_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_14_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_15_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_1_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_2_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_3_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_4_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_5_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_6_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_7_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_8_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_4_9_0_prog_clk));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout21 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net21));
 sky130_fd_sc_hd__buf_6 fanout22 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net23));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net25));
 sky130_fd_sc_hd__buf_6 fanout26 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out ),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_9_.out ),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out ),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_8_.out ),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out ),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_7_.out ),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out ),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_6_.out ),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out ),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_5_.out ),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out ),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_4_.out ),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out ),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_3_.out ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_2_.out ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_1_.out ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out ),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(\logical_tile_clb_mode_clb__0.mux_fle_0_in_0.INVTX1_0_.out ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_3_.Q ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_0_.Q ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_0_.Q ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_0_.Q ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_2_.Q ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_2_.Q ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_2_.Q ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_0_.Q ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_2_.Q ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_2_.Q ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_0_.Q ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_2_.Q ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_2_.Q ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_0_.Q ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_2_.Q ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_2_.Q ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_1_.Q ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_0_.Q ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_2_.Q ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_1_.Q ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_2_.Q ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_0_.Q ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_1_.Q ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_2_.Q ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_2_.Q ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_1_.Q ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_1_.Q ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_1_.Q ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_3.DFF_1_.Q ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_1_.Q ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_1_.Q ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_1_.Q ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_1_.Q ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_1_.Q ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_1_.Q ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_1_.Q ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_3_.Q ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_3_.Q ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_1_.Q ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.in ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.in ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.in ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.in ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.in ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.in ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.in ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.in ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.in ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_1.DFF_3_.Q ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.in ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.in ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.in ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.ccff_tail ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.in ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.in ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_2.DFF_3_.Q ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.DFF_0_.Q ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_1.DFF_3_.Q ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_3_.Q ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_3_.Q ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_3_.Q ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_0.DFF_3_.Q ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_3_.Q ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_3_.Q ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.in ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_2.DFF_0_.Q ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_0.DFF_0_.Q ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_3_.Q ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_3_.Q ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\logical_tile_clb_mode_clb__0.mem_fle_3_in_0.DFF_0_.Q ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_2.DFF_3_.Q ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_1.DFF_2_.Q ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_2_.Q ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_0_.Q ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_2.DFF_2_.Q ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_3.DFF_0_.Q ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\logical_tile_clb_mode_clb__0.mem_fle_1_in_0.DFF_0_.Q ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\logical_tile_clb_mode_clb__0.mem_fle_0_in_3.DFF_1_.Q ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_3.DFF_0_.Q ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\logical_tile_clb_mode_clb__0.mem_fle_2_in_1.DFF_0_.Q ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(bottom_width_0_height_0_subtile_0__pin_I_2_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(right_width_0_height_0_subtile_0__pin_I_9_),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(set),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(top_width_0_height_0_subtile_0__pin_I_0_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(top_width_0_height_0_subtile_0__pin_I_4_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(top_width_0_height_0_subtile_0__pin_I_8_),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input2 (.A(bottom_width_0_height_0_subtile_0__pin_I_6_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ccff_head),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(clk),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(left_width_0_height_0_subtile_0__pin_I_3_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(left_width_0_height_0_subtile_0__pin_I_7_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(reset),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(right_width_0_height_0_subtile_0__pin_I_1_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(right_width_0_height_0_subtile_0__pin_I_5_),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(bottom_width_0_height_0_subtile_0__pin_O_0_));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(ccff_tail));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(left_width_0_height_0_subtile_0__pin_O_1_));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(right_width_0_height_0_subtile_0__pin_O_3_));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(top_width_0_height_0_subtile_0__pin_O_2_));
endmodule

