magic
tech sky130A
magscale 1 2
timestamp 1708640337
<< viali >>
rect 15577 9605 15611 9639
rect 34253 9605 34287 9639
rect 36829 9605 36863 9639
rect 2053 9537 2087 9571
rect 4629 9537 4663 9571
rect 7205 9537 7239 9571
rect 9781 9537 9815 9571
rect 12357 9537 12391 9571
rect 18153 9537 18187 9571
rect 20729 9537 20763 9571
rect 23305 9537 23339 9571
rect 25881 9537 25915 9571
rect 29101 9537 29135 9571
rect 31677 9537 31711 9571
rect 38485 9537 38519 9571
rect 1409 9469 1443 9503
rect 38485 8857 38519 8891
rect 1409 8313 1443 8347
rect 38485 6205 38519 6239
rect 1409 5525 1443 5559
rect 38485 3485 38519 3519
rect 1409 2941 1443 2975
rect 13645 2397 13679 2431
rect 16221 2397 16255 2431
rect 18797 2397 18831 2431
rect 21373 2397 21407 2431
rect 23949 2397 23983 2431
rect 27169 2397 27203 2431
rect 37473 2397 37507 2431
rect 38485 2397 38519 2431
rect 1409 2261 1443 2295
rect 2697 2261 2731 2295
rect 5273 2261 5307 2295
rect 7849 2261 7883 2295
rect 10425 2261 10459 2295
rect 29745 2261 29779 2295
rect 32321 2261 32355 2295
rect 34897 2261 34931 2295
<< metal1 >>
rect 1104 9818 38984 9840
rect 1104 9766 10380 9818
rect 10432 9766 10444 9818
rect 10496 9766 10508 9818
rect 10560 9766 10572 9818
rect 10624 9766 10636 9818
rect 10688 9766 19810 9818
rect 19862 9766 19874 9818
rect 19926 9766 19938 9818
rect 19990 9766 20002 9818
rect 20054 9766 20066 9818
rect 20118 9766 29240 9818
rect 29292 9766 29304 9818
rect 29356 9766 29368 9818
rect 29420 9766 29432 9818
rect 29484 9766 29496 9818
rect 29548 9766 38670 9818
rect 38722 9766 38734 9818
rect 38786 9766 38798 9818
rect 38850 9766 38862 9818
rect 38914 9766 38926 9818
rect 38978 9766 38984 9818
rect 1104 9744 38984 9766
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 34238 9596 34244 9648
rect 34296 9596 34302 9648
rect 36814 9596 36820 9648
rect 36872 9596 36878 9648
rect 2038 9528 2044 9580
rect 2096 9528 2102 9580
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 18138 9528 18144 9580
rect 18196 9528 18202 9580
rect 20714 9528 20720 9580
rect 20772 9528 20778 9580
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 25866 9528 25872 9580
rect 25924 9528 25930 9580
rect 29086 9528 29092 9580
rect 29144 9528 29150 9580
rect 31662 9528 31668 9580
rect 31720 9528 31726 9580
rect 38470 9528 38476 9580
rect 38528 9528 38534 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2792 9500 2820 9528
rect 1443 9472 2820 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1104 9274 38824 9296
rect 1104 9222 5665 9274
rect 5717 9222 5729 9274
rect 5781 9222 5793 9274
rect 5845 9222 5857 9274
rect 5909 9222 5921 9274
rect 5973 9222 15095 9274
rect 15147 9222 15159 9274
rect 15211 9222 15223 9274
rect 15275 9222 15287 9274
rect 15339 9222 15351 9274
rect 15403 9222 24525 9274
rect 24577 9222 24589 9274
rect 24641 9222 24653 9274
rect 24705 9222 24717 9274
rect 24769 9222 24781 9274
rect 24833 9222 33955 9274
rect 34007 9222 34019 9274
rect 34071 9222 34083 9274
rect 34135 9222 34147 9274
rect 34199 9222 34211 9274
rect 34263 9222 38824 9274
rect 1104 9200 38824 9222
rect 38470 8848 38476 8900
rect 38528 8848 38534 8900
rect 1104 8730 38984 8752
rect 1104 8678 10380 8730
rect 10432 8678 10444 8730
rect 10496 8678 10508 8730
rect 10560 8678 10572 8730
rect 10624 8678 10636 8730
rect 10688 8678 19810 8730
rect 19862 8678 19874 8730
rect 19926 8678 19938 8730
rect 19990 8678 20002 8730
rect 20054 8678 20066 8730
rect 20118 8678 29240 8730
rect 29292 8678 29304 8730
rect 29356 8678 29368 8730
rect 29420 8678 29432 8730
rect 29484 8678 29496 8730
rect 29548 8678 38670 8730
rect 38722 8678 38734 8730
rect 38786 8678 38798 8730
rect 38850 8678 38862 8730
rect 38914 8678 38926 8730
rect 38978 8678 38984 8730
rect 1104 8656 38984 8678
rect 1394 8304 1400 8356
rect 1452 8304 1458 8356
rect 1104 8186 38824 8208
rect 1104 8134 5665 8186
rect 5717 8134 5729 8186
rect 5781 8134 5793 8186
rect 5845 8134 5857 8186
rect 5909 8134 5921 8186
rect 5973 8134 15095 8186
rect 15147 8134 15159 8186
rect 15211 8134 15223 8186
rect 15275 8134 15287 8186
rect 15339 8134 15351 8186
rect 15403 8134 24525 8186
rect 24577 8134 24589 8186
rect 24641 8134 24653 8186
rect 24705 8134 24717 8186
rect 24769 8134 24781 8186
rect 24833 8134 33955 8186
rect 34007 8134 34019 8186
rect 34071 8134 34083 8186
rect 34135 8134 34147 8186
rect 34199 8134 34211 8186
rect 34263 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38984 7664
rect 1104 7590 10380 7642
rect 10432 7590 10444 7642
rect 10496 7590 10508 7642
rect 10560 7590 10572 7642
rect 10624 7590 10636 7642
rect 10688 7590 19810 7642
rect 19862 7590 19874 7642
rect 19926 7590 19938 7642
rect 19990 7590 20002 7642
rect 20054 7590 20066 7642
rect 20118 7590 29240 7642
rect 29292 7590 29304 7642
rect 29356 7590 29368 7642
rect 29420 7590 29432 7642
rect 29484 7590 29496 7642
rect 29548 7590 38670 7642
rect 38722 7590 38734 7642
rect 38786 7590 38798 7642
rect 38850 7590 38862 7642
rect 38914 7590 38926 7642
rect 38978 7590 38984 7642
rect 1104 7568 38984 7590
rect 1104 7098 38824 7120
rect 1104 7046 5665 7098
rect 5717 7046 5729 7098
rect 5781 7046 5793 7098
rect 5845 7046 5857 7098
rect 5909 7046 5921 7098
rect 5973 7046 15095 7098
rect 15147 7046 15159 7098
rect 15211 7046 15223 7098
rect 15275 7046 15287 7098
rect 15339 7046 15351 7098
rect 15403 7046 24525 7098
rect 24577 7046 24589 7098
rect 24641 7046 24653 7098
rect 24705 7046 24717 7098
rect 24769 7046 24781 7098
rect 24833 7046 33955 7098
rect 34007 7046 34019 7098
rect 34071 7046 34083 7098
rect 34135 7046 34147 7098
rect 34199 7046 34211 7098
rect 34263 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38984 6576
rect 1104 6502 10380 6554
rect 10432 6502 10444 6554
rect 10496 6502 10508 6554
rect 10560 6502 10572 6554
rect 10624 6502 10636 6554
rect 10688 6502 19810 6554
rect 19862 6502 19874 6554
rect 19926 6502 19938 6554
rect 19990 6502 20002 6554
rect 20054 6502 20066 6554
rect 20118 6502 29240 6554
rect 29292 6502 29304 6554
rect 29356 6502 29368 6554
rect 29420 6502 29432 6554
rect 29484 6502 29496 6554
rect 29548 6502 38670 6554
rect 38722 6502 38734 6554
rect 38786 6502 38798 6554
rect 38850 6502 38862 6554
rect 38914 6502 38926 6554
rect 38978 6502 38984 6554
rect 1104 6480 38984 6502
rect 38470 6196 38476 6248
rect 38528 6196 38534 6248
rect 1104 6010 38824 6032
rect 1104 5958 5665 6010
rect 5717 5958 5729 6010
rect 5781 5958 5793 6010
rect 5845 5958 5857 6010
rect 5909 5958 5921 6010
rect 5973 5958 15095 6010
rect 15147 5958 15159 6010
rect 15211 5958 15223 6010
rect 15275 5958 15287 6010
rect 15339 5958 15351 6010
rect 15403 5958 24525 6010
rect 24577 5958 24589 6010
rect 24641 5958 24653 6010
rect 24705 5958 24717 6010
rect 24769 5958 24781 6010
rect 24833 5958 33955 6010
rect 34007 5958 34019 6010
rect 34071 5958 34083 6010
rect 34135 5958 34147 6010
rect 34199 5958 34211 6010
rect 34263 5958 38824 6010
rect 1104 5936 38824 5958
rect 1394 5516 1400 5568
rect 1452 5516 1458 5568
rect 1104 5466 38984 5488
rect 1104 5414 10380 5466
rect 10432 5414 10444 5466
rect 10496 5414 10508 5466
rect 10560 5414 10572 5466
rect 10624 5414 10636 5466
rect 10688 5414 19810 5466
rect 19862 5414 19874 5466
rect 19926 5414 19938 5466
rect 19990 5414 20002 5466
rect 20054 5414 20066 5466
rect 20118 5414 29240 5466
rect 29292 5414 29304 5466
rect 29356 5414 29368 5466
rect 29420 5414 29432 5466
rect 29484 5414 29496 5466
rect 29548 5414 38670 5466
rect 38722 5414 38734 5466
rect 38786 5414 38798 5466
rect 38850 5414 38862 5466
rect 38914 5414 38926 5466
rect 38978 5414 38984 5466
rect 1104 5392 38984 5414
rect 1104 4922 38824 4944
rect 1104 4870 5665 4922
rect 5717 4870 5729 4922
rect 5781 4870 5793 4922
rect 5845 4870 5857 4922
rect 5909 4870 5921 4922
rect 5973 4870 15095 4922
rect 15147 4870 15159 4922
rect 15211 4870 15223 4922
rect 15275 4870 15287 4922
rect 15339 4870 15351 4922
rect 15403 4870 24525 4922
rect 24577 4870 24589 4922
rect 24641 4870 24653 4922
rect 24705 4870 24717 4922
rect 24769 4870 24781 4922
rect 24833 4870 33955 4922
rect 34007 4870 34019 4922
rect 34071 4870 34083 4922
rect 34135 4870 34147 4922
rect 34199 4870 34211 4922
rect 34263 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38984 4400
rect 1104 4326 10380 4378
rect 10432 4326 10444 4378
rect 10496 4326 10508 4378
rect 10560 4326 10572 4378
rect 10624 4326 10636 4378
rect 10688 4326 19810 4378
rect 19862 4326 19874 4378
rect 19926 4326 19938 4378
rect 19990 4326 20002 4378
rect 20054 4326 20066 4378
rect 20118 4326 29240 4378
rect 29292 4326 29304 4378
rect 29356 4326 29368 4378
rect 29420 4326 29432 4378
rect 29484 4326 29496 4378
rect 29548 4326 38670 4378
rect 38722 4326 38734 4378
rect 38786 4326 38798 4378
rect 38850 4326 38862 4378
rect 38914 4326 38926 4378
rect 38978 4326 38984 4378
rect 1104 4304 38984 4326
rect 1104 3834 38824 3856
rect 1104 3782 5665 3834
rect 5717 3782 5729 3834
rect 5781 3782 5793 3834
rect 5845 3782 5857 3834
rect 5909 3782 5921 3834
rect 5973 3782 15095 3834
rect 15147 3782 15159 3834
rect 15211 3782 15223 3834
rect 15275 3782 15287 3834
rect 15339 3782 15351 3834
rect 15403 3782 24525 3834
rect 24577 3782 24589 3834
rect 24641 3782 24653 3834
rect 24705 3782 24717 3834
rect 24769 3782 24781 3834
rect 24833 3782 33955 3834
rect 34007 3782 34019 3834
rect 34071 3782 34083 3834
rect 34135 3782 34147 3834
rect 34199 3782 34211 3834
rect 34263 3782 38824 3834
rect 1104 3760 38824 3782
rect 38470 3476 38476 3528
rect 38528 3476 38534 3528
rect 1104 3290 38984 3312
rect 1104 3238 10380 3290
rect 10432 3238 10444 3290
rect 10496 3238 10508 3290
rect 10560 3238 10572 3290
rect 10624 3238 10636 3290
rect 10688 3238 19810 3290
rect 19862 3238 19874 3290
rect 19926 3238 19938 3290
rect 19990 3238 20002 3290
rect 20054 3238 20066 3290
rect 20118 3238 29240 3290
rect 29292 3238 29304 3290
rect 29356 3238 29368 3290
rect 29420 3238 29432 3290
rect 29484 3238 29496 3290
rect 29548 3238 38670 3290
rect 38722 3238 38734 3290
rect 38786 3238 38798 3290
rect 38850 3238 38862 3290
rect 38914 3238 38926 3290
rect 38978 3238 38984 3290
rect 1104 3216 38984 3238
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 992 2944 1409 2972
rect 992 2932 998 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1104 2746 38824 2768
rect 1104 2694 5665 2746
rect 5717 2694 5729 2746
rect 5781 2694 5793 2746
rect 5845 2694 5857 2746
rect 5909 2694 5921 2746
rect 5973 2694 15095 2746
rect 15147 2694 15159 2746
rect 15211 2694 15223 2746
rect 15275 2694 15287 2746
rect 15339 2694 15351 2746
rect 15403 2694 24525 2746
rect 24577 2694 24589 2746
rect 24641 2694 24653 2746
rect 24705 2694 24717 2746
rect 24769 2694 24781 2746
rect 24833 2694 33955 2746
rect 34007 2694 34019 2746
rect 34071 2694 34083 2746
rect 34135 2694 34147 2746
rect 34199 2694 34211 2746
rect 34263 2694 38824 2746
rect 1104 2672 38824 2694
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 21358 2388 21364 2440
rect 21416 2388 21422 2440
rect 23934 2388 23940 2440
rect 23992 2388 23998 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 290 2252 296 2304
rect 348 2292 354 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 348 2264 1409 2292
rect 348 2252 354 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 2682 2252 2688 2304
rect 2740 2252 2746 2304
rect 5258 2252 5264 2304
rect 5316 2252 5322 2304
rect 7834 2252 7840 2304
rect 7892 2252 7898 2304
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 10284 2264 10425 2292
rect 10284 2252 10290 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10413 2255 10471 2261
rect 29730 2252 29736 2304
rect 29788 2252 29794 2304
rect 32306 2252 32312 2304
rect 32364 2252 32370 2304
rect 34882 2252 34888 2304
rect 34940 2252 34946 2304
rect 1104 2202 38984 2224
rect 1104 2150 10380 2202
rect 10432 2150 10444 2202
rect 10496 2150 10508 2202
rect 10560 2150 10572 2202
rect 10624 2150 10636 2202
rect 10688 2150 19810 2202
rect 19862 2150 19874 2202
rect 19926 2150 19938 2202
rect 19990 2150 20002 2202
rect 20054 2150 20066 2202
rect 20118 2150 29240 2202
rect 29292 2150 29304 2202
rect 29356 2150 29368 2202
rect 29420 2150 29432 2202
rect 29484 2150 29496 2202
rect 29548 2150 38670 2202
rect 38722 2150 38734 2202
rect 38786 2150 38798 2202
rect 38850 2150 38862 2202
rect 38914 2150 38926 2202
rect 38978 2150 38984 2202
rect 1104 2128 38984 2150
<< via1 >>
rect 10380 9766 10432 9818
rect 10444 9766 10496 9818
rect 10508 9766 10560 9818
rect 10572 9766 10624 9818
rect 10636 9766 10688 9818
rect 19810 9766 19862 9818
rect 19874 9766 19926 9818
rect 19938 9766 19990 9818
rect 20002 9766 20054 9818
rect 20066 9766 20118 9818
rect 29240 9766 29292 9818
rect 29304 9766 29356 9818
rect 29368 9766 29420 9818
rect 29432 9766 29484 9818
rect 29496 9766 29548 9818
rect 38670 9766 38722 9818
rect 38734 9766 38786 9818
rect 38798 9766 38850 9818
rect 38862 9766 38914 9818
rect 38926 9766 38978 9818
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 34244 9639 34296 9648
rect 34244 9605 34253 9639
rect 34253 9605 34287 9639
rect 34287 9605 34296 9639
rect 34244 9596 34296 9605
rect 36820 9639 36872 9648
rect 36820 9605 36829 9639
rect 36829 9605 36863 9639
rect 36863 9605 36872 9639
rect 36820 9596 36872 9605
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2780 9528 2832 9580
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 25872 9571 25924 9580
rect 25872 9537 25881 9571
rect 25881 9537 25915 9571
rect 25915 9537 25924 9571
rect 25872 9528 25924 9537
rect 29092 9571 29144 9580
rect 29092 9537 29101 9571
rect 29101 9537 29135 9571
rect 29135 9537 29144 9571
rect 29092 9528 29144 9537
rect 31668 9571 31720 9580
rect 31668 9537 31677 9571
rect 31677 9537 31711 9571
rect 31711 9537 31720 9571
rect 31668 9528 31720 9537
rect 38476 9571 38528 9580
rect 38476 9537 38485 9571
rect 38485 9537 38519 9571
rect 38519 9537 38528 9571
rect 38476 9528 38528 9537
rect 5665 9222 5717 9274
rect 5729 9222 5781 9274
rect 5793 9222 5845 9274
rect 5857 9222 5909 9274
rect 5921 9222 5973 9274
rect 15095 9222 15147 9274
rect 15159 9222 15211 9274
rect 15223 9222 15275 9274
rect 15287 9222 15339 9274
rect 15351 9222 15403 9274
rect 24525 9222 24577 9274
rect 24589 9222 24641 9274
rect 24653 9222 24705 9274
rect 24717 9222 24769 9274
rect 24781 9222 24833 9274
rect 33955 9222 34007 9274
rect 34019 9222 34071 9274
rect 34083 9222 34135 9274
rect 34147 9222 34199 9274
rect 34211 9222 34263 9274
rect 38476 8891 38528 8900
rect 38476 8857 38485 8891
rect 38485 8857 38519 8891
rect 38519 8857 38528 8891
rect 38476 8848 38528 8857
rect 10380 8678 10432 8730
rect 10444 8678 10496 8730
rect 10508 8678 10560 8730
rect 10572 8678 10624 8730
rect 10636 8678 10688 8730
rect 19810 8678 19862 8730
rect 19874 8678 19926 8730
rect 19938 8678 19990 8730
rect 20002 8678 20054 8730
rect 20066 8678 20118 8730
rect 29240 8678 29292 8730
rect 29304 8678 29356 8730
rect 29368 8678 29420 8730
rect 29432 8678 29484 8730
rect 29496 8678 29548 8730
rect 38670 8678 38722 8730
rect 38734 8678 38786 8730
rect 38798 8678 38850 8730
rect 38862 8678 38914 8730
rect 38926 8678 38978 8730
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 5665 8134 5717 8186
rect 5729 8134 5781 8186
rect 5793 8134 5845 8186
rect 5857 8134 5909 8186
rect 5921 8134 5973 8186
rect 15095 8134 15147 8186
rect 15159 8134 15211 8186
rect 15223 8134 15275 8186
rect 15287 8134 15339 8186
rect 15351 8134 15403 8186
rect 24525 8134 24577 8186
rect 24589 8134 24641 8186
rect 24653 8134 24705 8186
rect 24717 8134 24769 8186
rect 24781 8134 24833 8186
rect 33955 8134 34007 8186
rect 34019 8134 34071 8186
rect 34083 8134 34135 8186
rect 34147 8134 34199 8186
rect 34211 8134 34263 8186
rect 10380 7590 10432 7642
rect 10444 7590 10496 7642
rect 10508 7590 10560 7642
rect 10572 7590 10624 7642
rect 10636 7590 10688 7642
rect 19810 7590 19862 7642
rect 19874 7590 19926 7642
rect 19938 7590 19990 7642
rect 20002 7590 20054 7642
rect 20066 7590 20118 7642
rect 29240 7590 29292 7642
rect 29304 7590 29356 7642
rect 29368 7590 29420 7642
rect 29432 7590 29484 7642
rect 29496 7590 29548 7642
rect 38670 7590 38722 7642
rect 38734 7590 38786 7642
rect 38798 7590 38850 7642
rect 38862 7590 38914 7642
rect 38926 7590 38978 7642
rect 5665 7046 5717 7098
rect 5729 7046 5781 7098
rect 5793 7046 5845 7098
rect 5857 7046 5909 7098
rect 5921 7046 5973 7098
rect 15095 7046 15147 7098
rect 15159 7046 15211 7098
rect 15223 7046 15275 7098
rect 15287 7046 15339 7098
rect 15351 7046 15403 7098
rect 24525 7046 24577 7098
rect 24589 7046 24641 7098
rect 24653 7046 24705 7098
rect 24717 7046 24769 7098
rect 24781 7046 24833 7098
rect 33955 7046 34007 7098
rect 34019 7046 34071 7098
rect 34083 7046 34135 7098
rect 34147 7046 34199 7098
rect 34211 7046 34263 7098
rect 10380 6502 10432 6554
rect 10444 6502 10496 6554
rect 10508 6502 10560 6554
rect 10572 6502 10624 6554
rect 10636 6502 10688 6554
rect 19810 6502 19862 6554
rect 19874 6502 19926 6554
rect 19938 6502 19990 6554
rect 20002 6502 20054 6554
rect 20066 6502 20118 6554
rect 29240 6502 29292 6554
rect 29304 6502 29356 6554
rect 29368 6502 29420 6554
rect 29432 6502 29484 6554
rect 29496 6502 29548 6554
rect 38670 6502 38722 6554
rect 38734 6502 38786 6554
rect 38798 6502 38850 6554
rect 38862 6502 38914 6554
rect 38926 6502 38978 6554
rect 38476 6239 38528 6248
rect 38476 6205 38485 6239
rect 38485 6205 38519 6239
rect 38519 6205 38528 6239
rect 38476 6196 38528 6205
rect 5665 5958 5717 6010
rect 5729 5958 5781 6010
rect 5793 5958 5845 6010
rect 5857 5958 5909 6010
rect 5921 5958 5973 6010
rect 15095 5958 15147 6010
rect 15159 5958 15211 6010
rect 15223 5958 15275 6010
rect 15287 5958 15339 6010
rect 15351 5958 15403 6010
rect 24525 5958 24577 6010
rect 24589 5958 24641 6010
rect 24653 5958 24705 6010
rect 24717 5958 24769 6010
rect 24781 5958 24833 6010
rect 33955 5958 34007 6010
rect 34019 5958 34071 6010
rect 34083 5958 34135 6010
rect 34147 5958 34199 6010
rect 34211 5958 34263 6010
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 10380 5414 10432 5466
rect 10444 5414 10496 5466
rect 10508 5414 10560 5466
rect 10572 5414 10624 5466
rect 10636 5414 10688 5466
rect 19810 5414 19862 5466
rect 19874 5414 19926 5466
rect 19938 5414 19990 5466
rect 20002 5414 20054 5466
rect 20066 5414 20118 5466
rect 29240 5414 29292 5466
rect 29304 5414 29356 5466
rect 29368 5414 29420 5466
rect 29432 5414 29484 5466
rect 29496 5414 29548 5466
rect 38670 5414 38722 5466
rect 38734 5414 38786 5466
rect 38798 5414 38850 5466
rect 38862 5414 38914 5466
rect 38926 5414 38978 5466
rect 5665 4870 5717 4922
rect 5729 4870 5781 4922
rect 5793 4870 5845 4922
rect 5857 4870 5909 4922
rect 5921 4870 5973 4922
rect 15095 4870 15147 4922
rect 15159 4870 15211 4922
rect 15223 4870 15275 4922
rect 15287 4870 15339 4922
rect 15351 4870 15403 4922
rect 24525 4870 24577 4922
rect 24589 4870 24641 4922
rect 24653 4870 24705 4922
rect 24717 4870 24769 4922
rect 24781 4870 24833 4922
rect 33955 4870 34007 4922
rect 34019 4870 34071 4922
rect 34083 4870 34135 4922
rect 34147 4870 34199 4922
rect 34211 4870 34263 4922
rect 10380 4326 10432 4378
rect 10444 4326 10496 4378
rect 10508 4326 10560 4378
rect 10572 4326 10624 4378
rect 10636 4326 10688 4378
rect 19810 4326 19862 4378
rect 19874 4326 19926 4378
rect 19938 4326 19990 4378
rect 20002 4326 20054 4378
rect 20066 4326 20118 4378
rect 29240 4326 29292 4378
rect 29304 4326 29356 4378
rect 29368 4326 29420 4378
rect 29432 4326 29484 4378
rect 29496 4326 29548 4378
rect 38670 4326 38722 4378
rect 38734 4326 38786 4378
rect 38798 4326 38850 4378
rect 38862 4326 38914 4378
rect 38926 4326 38978 4378
rect 5665 3782 5717 3834
rect 5729 3782 5781 3834
rect 5793 3782 5845 3834
rect 5857 3782 5909 3834
rect 5921 3782 5973 3834
rect 15095 3782 15147 3834
rect 15159 3782 15211 3834
rect 15223 3782 15275 3834
rect 15287 3782 15339 3834
rect 15351 3782 15403 3834
rect 24525 3782 24577 3834
rect 24589 3782 24641 3834
rect 24653 3782 24705 3834
rect 24717 3782 24769 3834
rect 24781 3782 24833 3834
rect 33955 3782 34007 3834
rect 34019 3782 34071 3834
rect 34083 3782 34135 3834
rect 34147 3782 34199 3834
rect 34211 3782 34263 3834
rect 38476 3519 38528 3528
rect 38476 3485 38485 3519
rect 38485 3485 38519 3519
rect 38519 3485 38528 3519
rect 38476 3476 38528 3485
rect 10380 3238 10432 3290
rect 10444 3238 10496 3290
rect 10508 3238 10560 3290
rect 10572 3238 10624 3290
rect 10636 3238 10688 3290
rect 19810 3238 19862 3290
rect 19874 3238 19926 3290
rect 19938 3238 19990 3290
rect 20002 3238 20054 3290
rect 20066 3238 20118 3290
rect 29240 3238 29292 3290
rect 29304 3238 29356 3290
rect 29368 3238 29420 3290
rect 29432 3238 29484 3290
rect 29496 3238 29548 3290
rect 38670 3238 38722 3290
rect 38734 3238 38786 3290
rect 38798 3238 38850 3290
rect 38862 3238 38914 3290
rect 38926 3238 38978 3290
rect 940 2932 992 2984
rect 5665 2694 5717 2746
rect 5729 2694 5781 2746
rect 5793 2694 5845 2746
rect 5857 2694 5909 2746
rect 5921 2694 5973 2746
rect 15095 2694 15147 2746
rect 15159 2694 15211 2746
rect 15223 2694 15275 2746
rect 15287 2694 15339 2746
rect 15351 2694 15403 2746
rect 24525 2694 24577 2746
rect 24589 2694 24641 2746
rect 24653 2694 24705 2746
rect 24717 2694 24769 2746
rect 24781 2694 24833 2746
rect 33955 2694 34007 2746
rect 34019 2694 34071 2746
rect 34083 2694 34135 2746
rect 34147 2694 34199 2746
rect 34211 2694 34263 2746
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 296 2252 348 2304
rect 2688 2295 2740 2304
rect 2688 2261 2697 2295
rect 2697 2261 2731 2295
rect 2731 2261 2740 2295
rect 2688 2252 2740 2261
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 7840 2295 7892 2304
rect 7840 2261 7849 2295
rect 7849 2261 7883 2295
rect 7883 2261 7892 2295
rect 7840 2252 7892 2261
rect 10232 2252 10284 2304
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 32312 2295 32364 2304
rect 32312 2261 32321 2295
rect 32321 2261 32355 2295
rect 32355 2261 32364 2295
rect 32312 2252 32364 2261
rect 34888 2295 34940 2304
rect 34888 2261 34897 2295
rect 34897 2261 34931 2295
rect 34931 2261 34940 2295
rect 34888 2252 34940 2261
rect 10380 2150 10432 2202
rect 10444 2150 10496 2202
rect 10508 2150 10560 2202
rect 10572 2150 10624 2202
rect 10636 2150 10688 2202
rect 19810 2150 19862 2202
rect 19874 2150 19926 2202
rect 19938 2150 19990 2202
rect 20002 2150 20054 2202
rect 20066 2150 20118 2202
rect 29240 2150 29292 2202
rect 29304 2150 29356 2202
rect 29368 2150 29420 2202
rect 29432 2150 29484 2202
rect 29496 2150 29548 2202
rect 38670 2150 38722 2202
rect 38734 2150 38786 2202
rect 38798 2150 38850 2202
rect 38862 2150 38914 2202
rect 38926 2150 38978 2202
<< metal2 >>
rect 1950 11200 2006 12000
rect 4526 11200 4582 12000
rect 7102 11200 7158 12000
rect 9678 11200 9734 12000
rect 12254 11200 12310 12000
rect 15474 11200 15530 12000
rect 18050 11200 18106 12000
rect 20626 11200 20682 12000
rect 23202 11200 23258 12000
rect 25778 11200 25834 12000
rect 28998 11200 29054 12000
rect 31574 11200 31630 12000
rect 34150 11200 34206 12000
rect 36726 11200 36782 12000
rect 38488 11206 39252 11234
rect 1964 9674 1992 11200
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 1964 9646 2084 9674
rect 2056 9586 2084 9646
rect 2792 9586 2820 10911
rect 4540 9674 4568 11200
rect 7116 9674 7144 11200
rect 9692 9674 9720 11200
rect 10380 9820 10688 9829
rect 10380 9818 10386 9820
rect 10442 9818 10466 9820
rect 10522 9818 10546 9820
rect 10602 9818 10626 9820
rect 10682 9818 10688 9820
rect 10442 9766 10444 9818
rect 10624 9766 10626 9818
rect 10380 9764 10386 9766
rect 10442 9764 10466 9766
rect 10522 9764 10546 9766
rect 10602 9764 10626 9766
rect 10682 9764 10688 9766
rect 10380 9755 10688 9764
rect 12268 9674 12296 11200
rect 15488 9674 15516 11200
rect 18064 9674 18092 11200
rect 19810 9820 20118 9829
rect 19810 9818 19816 9820
rect 19872 9818 19896 9820
rect 19952 9818 19976 9820
rect 20032 9818 20056 9820
rect 20112 9818 20118 9820
rect 19872 9766 19874 9818
rect 20054 9766 20056 9818
rect 19810 9764 19816 9766
rect 19872 9764 19896 9766
rect 19952 9764 19976 9766
rect 20032 9764 20056 9766
rect 20112 9764 20118 9766
rect 19810 9755 20118 9764
rect 20640 9674 20668 11200
rect 23216 9674 23244 11200
rect 25792 9674 25820 11200
rect 29012 9674 29040 11200
rect 29240 9820 29548 9829
rect 29240 9818 29246 9820
rect 29302 9818 29326 9820
rect 29382 9818 29406 9820
rect 29462 9818 29486 9820
rect 29542 9818 29548 9820
rect 29302 9766 29304 9818
rect 29484 9766 29486 9818
rect 29240 9764 29246 9766
rect 29302 9764 29326 9766
rect 29382 9764 29406 9766
rect 29462 9764 29486 9766
rect 29542 9764 29548 9766
rect 29240 9755 29548 9764
rect 31588 9674 31616 11200
rect 34164 9674 34192 11200
rect 36740 9674 36768 11200
rect 4540 9646 4660 9674
rect 7116 9646 7236 9674
rect 9692 9646 9812 9674
rect 12268 9646 12388 9674
rect 15488 9654 15608 9674
rect 15488 9648 15620 9654
rect 15488 9646 15568 9648
rect 4632 9586 4660 9646
rect 7208 9586 7236 9646
rect 9784 9586 9812 9646
rect 12360 9586 12388 9646
rect 18064 9646 18184 9674
rect 20640 9646 20760 9674
rect 23216 9646 23336 9674
rect 25792 9646 25912 9674
rect 29012 9646 29132 9674
rect 31588 9646 31708 9674
rect 34164 9654 34284 9674
rect 36740 9654 36860 9674
rect 34164 9648 34296 9654
rect 34164 9646 34244 9648
rect 15568 9590 15620 9596
rect 18156 9586 18184 9646
rect 20732 9586 20760 9646
rect 23308 9586 23336 9646
rect 25884 9586 25912 9646
rect 29104 9586 29132 9646
rect 31680 9586 31708 9646
rect 36740 9648 36872 9654
rect 36740 9646 36820 9648
rect 34244 9590 34296 9596
rect 36820 9590 36872 9596
rect 38488 9586 38516 11206
rect 39224 11098 39252 11206
rect 39302 11200 39358 12000
rect 39316 11098 39344 11200
rect 39224 11070 39344 11098
rect 38670 9820 38978 9829
rect 38670 9818 38676 9820
rect 38732 9818 38756 9820
rect 38812 9818 38836 9820
rect 38892 9818 38916 9820
rect 38972 9818 38978 9820
rect 38732 9766 38734 9818
rect 38914 9766 38916 9818
rect 38670 9764 38676 9766
rect 38732 9764 38756 9766
rect 38812 9764 38836 9766
rect 38892 9764 38916 9766
rect 38972 9764 38978 9766
rect 38670 9755 38978 9764
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 38476 9580 38528 9586
rect 38476 9522 38528 9528
rect 5665 9276 5973 9285
rect 5665 9274 5671 9276
rect 5727 9274 5751 9276
rect 5807 9274 5831 9276
rect 5887 9274 5911 9276
rect 5967 9274 5973 9276
rect 5727 9222 5729 9274
rect 5909 9222 5911 9274
rect 5665 9220 5671 9222
rect 5727 9220 5751 9222
rect 5807 9220 5831 9222
rect 5887 9220 5911 9222
rect 5967 9220 5973 9222
rect 5665 9211 5973 9220
rect 15095 9276 15403 9285
rect 15095 9274 15101 9276
rect 15157 9274 15181 9276
rect 15237 9274 15261 9276
rect 15317 9274 15341 9276
rect 15397 9274 15403 9276
rect 15157 9222 15159 9274
rect 15339 9222 15341 9274
rect 15095 9220 15101 9222
rect 15157 9220 15181 9222
rect 15237 9220 15261 9222
rect 15317 9220 15341 9222
rect 15397 9220 15403 9222
rect 15095 9211 15403 9220
rect 24525 9276 24833 9285
rect 24525 9274 24531 9276
rect 24587 9274 24611 9276
rect 24667 9274 24691 9276
rect 24747 9274 24771 9276
rect 24827 9274 24833 9276
rect 24587 9222 24589 9274
rect 24769 9222 24771 9274
rect 24525 9220 24531 9222
rect 24587 9220 24611 9222
rect 24667 9220 24691 9222
rect 24747 9220 24771 9222
rect 24827 9220 24833 9222
rect 24525 9211 24833 9220
rect 33955 9276 34263 9285
rect 33955 9274 33961 9276
rect 34017 9274 34041 9276
rect 34097 9274 34121 9276
rect 34177 9274 34201 9276
rect 34257 9274 34263 9276
rect 34017 9222 34019 9274
rect 34199 9222 34201 9274
rect 33955 9220 33961 9222
rect 34017 9220 34041 9222
rect 34097 9220 34121 9222
rect 34177 9220 34201 9222
rect 34257 9220 34263 9222
rect 33955 9211 34263 9220
rect 38474 8936 38530 8945
rect 38474 8871 38476 8880
rect 38528 8871 38530 8880
rect 38476 8842 38528 8848
rect 10380 8732 10688 8741
rect 10380 8730 10386 8732
rect 10442 8730 10466 8732
rect 10522 8730 10546 8732
rect 10602 8730 10626 8732
rect 10682 8730 10688 8732
rect 10442 8678 10444 8730
rect 10624 8678 10626 8730
rect 10380 8676 10386 8678
rect 10442 8676 10466 8678
rect 10522 8676 10546 8678
rect 10602 8676 10626 8678
rect 10682 8676 10688 8678
rect 10380 8667 10688 8676
rect 19810 8732 20118 8741
rect 19810 8730 19816 8732
rect 19872 8730 19896 8732
rect 19952 8730 19976 8732
rect 20032 8730 20056 8732
rect 20112 8730 20118 8732
rect 19872 8678 19874 8730
rect 20054 8678 20056 8730
rect 19810 8676 19816 8678
rect 19872 8676 19896 8678
rect 19952 8676 19976 8678
rect 20032 8676 20056 8678
rect 20112 8676 20118 8678
rect 19810 8667 20118 8676
rect 29240 8732 29548 8741
rect 29240 8730 29246 8732
rect 29302 8730 29326 8732
rect 29382 8730 29406 8732
rect 29462 8730 29486 8732
rect 29542 8730 29548 8732
rect 29302 8678 29304 8730
rect 29484 8678 29486 8730
rect 29240 8676 29246 8678
rect 29302 8676 29326 8678
rect 29382 8676 29406 8678
rect 29462 8676 29486 8678
rect 29542 8676 29548 8678
rect 29240 8667 29548 8676
rect 38670 8732 38978 8741
rect 38670 8730 38676 8732
rect 38732 8730 38756 8732
rect 38812 8730 38836 8732
rect 38892 8730 38916 8732
rect 38972 8730 38978 8732
rect 38732 8678 38734 8730
rect 38914 8678 38916 8730
rect 38670 8676 38676 8678
rect 38732 8676 38756 8678
rect 38812 8676 38836 8678
rect 38892 8676 38916 8678
rect 38972 8676 38978 8678
rect 38670 8667 38978 8676
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 5665 8188 5973 8197
rect 5665 8186 5671 8188
rect 5727 8186 5751 8188
rect 5807 8186 5831 8188
rect 5887 8186 5911 8188
rect 5967 8186 5973 8188
rect 5727 8134 5729 8186
rect 5909 8134 5911 8186
rect 5665 8132 5671 8134
rect 5727 8132 5751 8134
rect 5807 8132 5831 8134
rect 5887 8132 5911 8134
rect 5967 8132 5973 8134
rect 5665 8123 5973 8132
rect 15095 8188 15403 8197
rect 15095 8186 15101 8188
rect 15157 8186 15181 8188
rect 15237 8186 15261 8188
rect 15317 8186 15341 8188
rect 15397 8186 15403 8188
rect 15157 8134 15159 8186
rect 15339 8134 15341 8186
rect 15095 8132 15101 8134
rect 15157 8132 15181 8134
rect 15237 8132 15261 8134
rect 15317 8132 15341 8134
rect 15397 8132 15403 8134
rect 15095 8123 15403 8132
rect 24525 8188 24833 8197
rect 24525 8186 24531 8188
rect 24587 8186 24611 8188
rect 24667 8186 24691 8188
rect 24747 8186 24771 8188
rect 24827 8186 24833 8188
rect 24587 8134 24589 8186
rect 24769 8134 24771 8186
rect 24525 8132 24531 8134
rect 24587 8132 24611 8134
rect 24667 8132 24691 8134
rect 24747 8132 24771 8134
rect 24827 8132 24833 8134
rect 24525 8123 24833 8132
rect 33955 8188 34263 8197
rect 33955 8186 33961 8188
rect 34017 8186 34041 8188
rect 34097 8186 34121 8188
rect 34177 8186 34201 8188
rect 34257 8186 34263 8188
rect 34017 8134 34019 8186
rect 34199 8134 34201 8186
rect 33955 8132 33961 8134
rect 34017 8132 34041 8134
rect 34097 8132 34121 8134
rect 34177 8132 34201 8134
rect 34257 8132 34263 8134
rect 33955 8123 34263 8132
rect 10380 7644 10688 7653
rect 10380 7642 10386 7644
rect 10442 7642 10466 7644
rect 10522 7642 10546 7644
rect 10602 7642 10626 7644
rect 10682 7642 10688 7644
rect 10442 7590 10444 7642
rect 10624 7590 10626 7642
rect 10380 7588 10386 7590
rect 10442 7588 10466 7590
rect 10522 7588 10546 7590
rect 10602 7588 10626 7590
rect 10682 7588 10688 7590
rect 10380 7579 10688 7588
rect 19810 7644 20118 7653
rect 19810 7642 19816 7644
rect 19872 7642 19896 7644
rect 19952 7642 19976 7644
rect 20032 7642 20056 7644
rect 20112 7642 20118 7644
rect 19872 7590 19874 7642
rect 20054 7590 20056 7642
rect 19810 7588 19816 7590
rect 19872 7588 19896 7590
rect 19952 7588 19976 7590
rect 20032 7588 20056 7590
rect 20112 7588 20118 7590
rect 19810 7579 20118 7588
rect 29240 7644 29548 7653
rect 29240 7642 29246 7644
rect 29302 7642 29326 7644
rect 29382 7642 29406 7644
rect 29462 7642 29486 7644
rect 29542 7642 29548 7644
rect 29302 7590 29304 7642
rect 29484 7590 29486 7642
rect 29240 7588 29246 7590
rect 29302 7588 29326 7590
rect 29382 7588 29406 7590
rect 29462 7588 29486 7590
rect 29542 7588 29548 7590
rect 29240 7579 29548 7588
rect 38670 7644 38978 7653
rect 38670 7642 38676 7644
rect 38732 7642 38756 7644
rect 38812 7642 38836 7644
rect 38892 7642 38916 7644
rect 38972 7642 38978 7644
rect 38732 7590 38734 7642
rect 38914 7590 38916 7642
rect 38670 7588 38676 7590
rect 38732 7588 38756 7590
rect 38812 7588 38836 7590
rect 38892 7588 38916 7590
rect 38972 7588 38978 7590
rect 38670 7579 38978 7588
rect 5665 7100 5973 7109
rect 5665 7098 5671 7100
rect 5727 7098 5751 7100
rect 5807 7098 5831 7100
rect 5887 7098 5911 7100
rect 5967 7098 5973 7100
rect 5727 7046 5729 7098
rect 5909 7046 5911 7098
rect 5665 7044 5671 7046
rect 5727 7044 5751 7046
rect 5807 7044 5831 7046
rect 5887 7044 5911 7046
rect 5967 7044 5973 7046
rect 5665 7035 5973 7044
rect 15095 7100 15403 7109
rect 15095 7098 15101 7100
rect 15157 7098 15181 7100
rect 15237 7098 15261 7100
rect 15317 7098 15341 7100
rect 15397 7098 15403 7100
rect 15157 7046 15159 7098
rect 15339 7046 15341 7098
rect 15095 7044 15101 7046
rect 15157 7044 15181 7046
rect 15237 7044 15261 7046
rect 15317 7044 15341 7046
rect 15397 7044 15403 7046
rect 15095 7035 15403 7044
rect 24525 7100 24833 7109
rect 24525 7098 24531 7100
rect 24587 7098 24611 7100
rect 24667 7098 24691 7100
rect 24747 7098 24771 7100
rect 24827 7098 24833 7100
rect 24587 7046 24589 7098
rect 24769 7046 24771 7098
rect 24525 7044 24531 7046
rect 24587 7044 24611 7046
rect 24667 7044 24691 7046
rect 24747 7044 24771 7046
rect 24827 7044 24833 7046
rect 24525 7035 24833 7044
rect 33955 7100 34263 7109
rect 33955 7098 33961 7100
rect 34017 7098 34041 7100
rect 34097 7098 34121 7100
rect 34177 7098 34201 7100
rect 34257 7098 34263 7100
rect 34017 7046 34019 7098
rect 34199 7046 34201 7098
rect 33955 7044 33961 7046
rect 34017 7044 34041 7046
rect 34097 7044 34121 7046
rect 34177 7044 34201 7046
rect 34257 7044 34263 7046
rect 33955 7035 34263 7044
rect 10380 6556 10688 6565
rect 10380 6554 10386 6556
rect 10442 6554 10466 6556
rect 10522 6554 10546 6556
rect 10602 6554 10626 6556
rect 10682 6554 10688 6556
rect 10442 6502 10444 6554
rect 10624 6502 10626 6554
rect 10380 6500 10386 6502
rect 10442 6500 10466 6502
rect 10522 6500 10546 6502
rect 10602 6500 10626 6502
rect 10682 6500 10688 6502
rect 10380 6491 10688 6500
rect 19810 6556 20118 6565
rect 19810 6554 19816 6556
rect 19872 6554 19896 6556
rect 19952 6554 19976 6556
rect 20032 6554 20056 6556
rect 20112 6554 20118 6556
rect 19872 6502 19874 6554
rect 20054 6502 20056 6554
rect 19810 6500 19816 6502
rect 19872 6500 19896 6502
rect 19952 6500 19976 6502
rect 20032 6500 20056 6502
rect 20112 6500 20118 6502
rect 19810 6491 20118 6500
rect 29240 6556 29548 6565
rect 29240 6554 29246 6556
rect 29302 6554 29326 6556
rect 29382 6554 29406 6556
rect 29462 6554 29486 6556
rect 29542 6554 29548 6556
rect 29302 6502 29304 6554
rect 29484 6502 29486 6554
rect 29240 6500 29246 6502
rect 29302 6500 29326 6502
rect 29382 6500 29406 6502
rect 29462 6500 29486 6502
rect 29542 6500 29548 6502
rect 29240 6491 29548 6500
rect 38670 6556 38978 6565
rect 38670 6554 38676 6556
rect 38732 6554 38756 6556
rect 38812 6554 38836 6556
rect 38892 6554 38916 6556
rect 38972 6554 38978 6556
rect 38732 6502 38734 6554
rect 38914 6502 38916 6554
rect 38670 6500 38676 6502
rect 38732 6500 38756 6502
rect 38812 6500 38836 6502
rect 38892 6500 38916 6502
rect 38972 6500 38978 6502
rect 38670 6491 38978 6500
rect 38476 6248 38528 6254
rect 38474 6216 38476 6225
rect 38528 6216 38530 6225
rect 38474 6151 38530 6160
rect 5665 6012 5973 6021
rect 5665 6010 5671 6012
rect 5727 6010 5751 6012
rect 5807 6010 5831 6012
rect 5887 6010 5911 6012
rect 5967 6010 5973 6012
rect 5727 5958 5729 6010
rect 5909 5958 5911 6010
rect 5665 5956 5671 5958
rect 5727 5956 5751 5958
rect 5807 5956 5831 5958
rect 5887 5956 5911 5958
rect 5967 5956 5973 5958
rect 5665 5947 5973 5956
rect 15095 6012 15403 6021
rect 15095 6010 15101 6012
rect 15157 6010 15181 6012
rect 15237 6010 15261 6012
rect 15317 6010 15341 6012
rect 15397 6010 15403 6012
rect 15157 5958 15159 6010
rect 15339 5958 15341 6010
rect 15095 5956 15101 5958
rect 15157 5956 15181 5958
rect 15237 5956 15261 5958
rect 15317 5956 15341 5958
rect 15397 5956 15403 5958
rect 15095 5947 15403 5956
rect 24525 6012 24833 6021
rect 24525 6010 24531 6012
rect 24587 6010 24611 6012
rect 24667 6010 24691 6012
rect 24747 6010 24771 6012
rect 24827 6010 24833 6012
rect 24587 5958 24589 6010
rect 24769 5958 24771 6010
rect 24525 5956 24531 5958
rect 24587 5956 24611 5958
rect 24667 5956 24691 5958
rect 24747 5956 24771 5958
rect 24827 5956 24833 5958
rect 24525 5947 24833 5956
rect 33955 6012 34263 6021
rect 33955 6010 33961 6012
rect 34017 6010 34041 6012
rect 34097 6010 34121 6012
rect 34177 6010 34201 6012
rect 34257 6010 34263 6012
rect 34017 5958 34019 6010
rect 34199 5958 34201 6010
rect 33955 5956 33961 5958
rect 34017 5956 34041 5958
rect 34097 5956 34121 5958
rect 34177 5956 34201 5958
rect 34257 5956 34263 5958
rect 33955 5947 34263 5956
rect 1400 5568 1452 5574
rect 1398 5536 1400 5545
rect 1452 5536 1454 5545
rect 1398 5471 1454 5480
rect 10380 5468 10688 5477
rect 10380 5466 10386 5468
rect 10442 5466 10466 5468
rect 10522 5466 10546 5468
rect 10602 5466 10626 5468
rect 10682 5466 10688 5468
rect 10442 5414 10444 5466
rect 10624 5414 10626 5466
rect 10380 5412 10386 5414
rect 10442 5412 10466 5414
rect 10522 5412 10546 5414
rect 10602 5412 10626 5414
rect 10682 5412 10688 5414
rect 10380 5403 10688 5412
rect 19810 5468 20118 5477
rect 19810 5466 19816 5468
rect 19872 5466 19896 5468
rect 19952 5466 19976 5468
rect 20032 5466 20056 5468
rect 20112 5466 20118 5468
rect 19872 5414 19874 5466
rect 20054 5414 20056 5466
rect 19810 5412 19816 5414
rect 19872 5412 19896 5414
rect 19952 5412 19976 5414
rect 20032 5412 20056 5414
rect 20112 5412 20118 5414
rect 19810 5403 20118 5412
rect 29240 5468 29548 5477
rect 29240 5466 29246 5468
rect 29302 5466 29326 5468
rect 29382 5466 29406 5468
rect 29462 5466 29486 5468
rect 29542 5466 29548 5468
rect 29302 5414 29304 5466
rect 29484 5414 29486 5466
rect 29240 5412 29246 5414
rect 29302 5412 29326 5414
rect 29382 5412 29406 5414
rect 29462 5412 29486 5414
rect 29542 5412 29548 5414
rect 29240 5403 29548 5412
rect 38670 5468 38978 5477
rect 38670 5466 38676 5468
rect 38732 5466 38756 5468
rect 38812 5466 38836 5468
rect 38892 5466 38916 5468
rect 38972 5466 38978 5468
rect 38732 5414 38734 5466
rect 38914 5414 38916 5466
rect 38670 5412 38676 5414
rect 38732 5412 38756 5414
rect 38812 5412 38836 5414
rect 38892 5412 38916 5414
rect 38972 5412 38978 5414
rect 38670 5403 38978 5412
rect 5665 4924 5973 4933
rect 5665 4922 5671 4924
rect 5727 4922 5751 4924
rect 5807 4922 5831 4924
rect 5887 4922 5911 4924
rect 5967 4922 5973 4924
rect 5727 4870 5729 4922
rect 5909 4870 5911 4922
rect 5665 4868 5671 4870
rect 5727 4868 5751 4870
rect 5807 4868 5831 4870
rect 5887 4868 5911 4870
rect 5967 4868 5973 4870
rect 5665 4859 5973 4868
rect 15095 4924 15403 4933
rect 15095 4922 15101 4924
rect 15157 4922 15181 4924
rect 15237 4922 15261 4924
rect 15317 4922 15341 4924
rect 15397 4922 15403 4924
rect 15157 4870 15159 4922
rect 15339 4870 15341 4922
rect 15095 4868 15101 4870
rect 15157 4868 15181 4870
rect 15237 4868 15261 4870
rect 15317 4868 15341 4870
rect 15397 4868 15403 4870
rect 15095 4859 15403 4868
rect 24525 4924 24833 4933
rect 24525 4922 24531 4924
rect 24587 4922 24611 4924
rect 24667 4922 24691 4924
rect 24747 4922 24771 4924
rect 24827 4922 24833 4924
rect 24587 4870 24589 4922
rect 24769 4870 24771 4922
rect 24525 4868 24531 4870
rect 24587 4868 24611 4870
rect 24667 4868 24691 4870
rect 24747 4868 24771 4870
rect 24827 4868 24833 4870
rect 24525 4859 24833 4868
rect 33955 4924 34263 4933
rect 33955 4922 33961 4924
rect 34017 4922 34041 4924
rect 34097 4922 34121 4924
rect 34177 4922 34201 4924
rect 34257 4922 34263 4924
rect 34017 4870 34019 4922
rect 34199 4870 34201 4922
rect 33955 4868 33961 4870
rect 34017 4868 34041 4870
rect 34097 4868 34121 4870
rect 34177 4868 34201 4870
rect 34257 4868 34263 4870
rect 33955 4859 34263 4868
rect 10380 4380 10688 4389
rect 10380 4378 10386 4380
rect 10442 4378 10466 4380
rect 10522 4378 10546 4380
rect 10602 4378 10626 4380
rect 10682 4378 10688 4380
rect 10442 4326 10444 4378
rect 10624 4326 10626 4378
rect 10380 4324 10386 4326
rect 10442 4324 10466 4326
rect 10522 4324 10546 4326
rect 10602 4324 10626 4326
rect 10682 4324 10688 4326
rect 10380 4315 10688 4324
rect 19810 4380 20118 4389
rect 19810 4378 19816 4380
rect 19872 4378 19896 4380
rect 19952 4378 19976 4380
rect 20032 4378 20056 4380
rect 20112 4378 20118 4380
rect 19872 4326 19874 4378
rect 20054 4326 20056 4378
rect 19810 4324 19816 4326
rect 19872 4324 19896 4326
rect 19952 4324 19976 4326
rect 20032 4324 20056 4326
rect 20112 4324 20118 4326
rect 19810 4315 20118 4324
rect 29240 4380 29548 4389
rect 29240 4378 29246 4380
rect 29302 4378 29326 4380
rect 29382 4378 29406 4380
rect 29462 4378 29486 4380
rect 29542 4378 29548 4380
rect 29302 4326 29304 4378
rect 29484 4326 29486 4378
rect 29240 4324 29246 4326
rect 29302 4324 29326 4326
rect 29382 4324 29406 4326
rect 29462 4324 29486 4326
rect 29542 4324 29548 4326
rect 29240 4315 29548 4324
rect 38670 4380 38978 4389
rect 38670 4378 38676 4380
rect 38732 4378 38756 4380
rect 38812 4378 38836 4380
rect 38892 4378 38916 4380
rect 38972 4378 38978 4380
rect 38732 4326 38734 4378
rect 38914 4326 38916 4378
rect 38670 4324 38676 4326
rect 38732 4324 38756 4326
rect 38812 4324 38836 4326
rect 38892 4324 38916 4326
rect 38972 4324 38978 4326
rect 38670 4315 38978 4324
rect 5665 3836 5973 3845
rect 5665 3834 5671 3836
rect 5727 3834 5751 3836
rect 5807 3834 5831 3836
rect 5887 3834 5911 3836
rect 5967 3834 5973 3836
rect 5727 3782 5729 3834
rect 5909 3782 5911 3834
rect 5665 3780 5671 3782
rect 5727 3780 5751 3782
rect 5807 3780 5831 3782
rect 5887 3780 5911 3782
rect 5967 3780 5973 3782
rect 5665 3771 5973 3780
rect 15095 3836 15403 3845
rect 15095 3834 15101 3836
rect 15157 3834 15181 3836
rect 15237 3834 15261 3836
rect 15317 3834 15341 3836
rect 15397 3834 15403 3836
rect 15157 3782 15159 3834
rect 15339 3782 15341 3834
rect 15095 3780 15101 3782
rect 15157 3780 15181 3782
rect 15237 3780 15261 3782
rect 15317 3780 15341 3782
rect 15397 3780 15403 3782
rect 15095 3771 15403 3780
rect 24525 3836 24833 3845
rect 24525 3834 24531 3836
rect 24587 3834 24611 3836
rect 24667 3834 24691 3836
rect 24747 3834 24771 3836
rect 24827 3834 24833 3836
rect 24587 3782 24589 3834
rect 24769 3782 24771 3834
rect 24525 3780 24531 3782
rect 24587 3780 24611 3782
rect 24667 3780 24691 3782
rect 24747 3780 24771 3782
rect 24827 3780 24833 3782
rect 24525 3771 24833 3780
rect 33955 3836 34263 3845
rect 33955 3834 33961 3836
rect 34017 3834 34041 3836
rect 34097 3834 34121 3836
rect 34177 3834 34201 3836
rect 34257 3834 34263 3836
rect 34017 3782 34019 3834
rect 34199 3782 34201 3834
rect 33955 3780 33961 3782
rect 34017 3780 34041 3782
rect 34097 3780 34121 3782
rect 34177 3780 34201 3782
rect 34257 3780 34263 3782
rect 33955 3771 34263 3780
rect 38476 3528 38528 3534
rect 38474 3496 38476 3505
rect 38528 3496 38530 3505
rect 38474 3431 38530 3440
rect 10380 3292 10688 3301
rect 10380 3290 10386 3292
rect 10442 3290 10466 3292
rect 10522 3290 10546 3292
rect 10602 3290 10626 3292
rect 10682 3290 10688 3292
rect 10442 3238 10444 3290
rect 10624 3238 10626 3290
rect 10380 3236 10386 3238
rect 10442 3236 10466 3238
rect 10522 3236 10546 3238
rect 10602 3236 10626 3238
rect 10682 3236 10688 3238
rect 10380 3227 10688 3236
rect 19810 3292 20118 3301
rect 19810 3290 19816 3292
rect 19872 3290 19896 3292
rect 19952 3290 19976 3292
rect 20032 3290 20056 3292
rect 20112 3290 20118 3292
rect 19872 3238 19874 3290
rect 20054 3238 20056 3290
rect 19810 3236 19816 3238
rect 19872 3236 19896 3238
rect 19952 3236 19976 3238
rect 20032 3236 20056 3238
rect 20112 3236 20118 3238
rect 19810 3227 20118 3236
rect 29240 3292 29548 3301
rect 29240 3290 29246 3292
rect 29302 3290 29326 3292
rect 29382 3290 29406 3292
rect 29462 3290 29486 3292
rect 29542 3290 29548 3292
rect 29302 3238 29304 3290
rect 29484 3238 29486 3290
rect 29240 3236 29246 3238
rect 29302 3236 29326 3238
rect 29382 3236 29406 3238
rect 29462 3236 29486 3238
rect 29542 3236 29548 3238
rect 29240 3227 29548 3236
rect 38670 3292 38978 3301
rect 38670 3290 38676 3292
rect 38732 3290 38756 3292
rect 38812 3290 38836 3292
rect 38892 3290 38916 3292
rect 38972 3290 38978 3292
rect 38732 3238 38734 3290
rect 38914 3238 38916 3290
rect 38670 3236 38676 3238
rect 38732 3236 38756 3238
rect 38812 3236 38836 3238
rect 38892 3236 38916 3238
rect 38972 3236 38978 3238
rect 38670 3227 38978 3236
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 2825 980 2926
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 5665 2748 5973 2757
rect 5665 2746 5671 2748
rect 5727 2746 5751 2748
rect 5807 2746 5831 2748
rect 5887 2746 5911 2748
rect 5967 2746 5973 2748
rect 5727 2694 5729 2746
rect 5909 2694 5911 2746
rect 5665 2692 5671 2694
rect 5727 2692 5751 2694
rect 5807 2692 5831 2694
rect 5887 2692 5911 2694
rect 5967 2692 5973 2694
rect 5665 2683 5973 2692
rect 15095 2748 15403 2757
rect 15095 2746 15101 2748
rect 15157 2746 15181 2748
rect 15237 2746 15261 2748
rect 15317 2746 15341 2748
rect 15397 2746 15403 2748
rect 15157 2694 15159 2746
rect 15339 2694 15341 2746
rect 15095 2692 15101 2694
rect 15157 2692 15181 2694
rect 15237 2692 15261 2694
rect 15317 2692 15341 2694
rect 15397 2692 15403 2694
rect 15095 2683 15403 2692
rect 24525 2748 24833 2757
rect 24525 2746 24531 2748
rect 24587 2746 24611 2748
rect 24667 2746 24691 2748
rect 24747 2746 24771 2748
rect 24827 2746 24833 2748
rect 24587 2694 24589 2746
rect 24769 2694 24771 2746
rect 24525 2692 24531 2694
rect 24587 2692 24611 2694
rect 24667 2692 24691 2694
rect 24747 2692 24771 2694
rect 24827 2692 24833 2694
rect 24525 2683 24833 2692
rect 33955 2748 34263 2757
rect 33955 2746 33961 2748
rect 34017 2746 34041 2748
rect 34097 2746 34121 2748
rect 34177 2746 34201 2748
rect 34257 2746 34263 2748
rect 34017 2694 34019 2746
rect 34199 2694 34201 2746
rect 33955 2692 33961 2694
rect 34017 2692 34041 2694
rect 34097 2692 34121 2694
rect 34177 2692 34201 2694
rect 34257 2692 34263 2694
rect 33955 2683 34263 2692
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 296 2304 348 2310
rect 296 2246 348 2252
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 32 870 152 898
rect 32 800 60 870
rect 18 0 74 800
rect 124 762 152 870
rect 308 762 336 2246
rect 2700 1170 2728 2246
rect 5276 1170 5304 2246
rect 7852 1170 7880 2246
rect 2608 1142 2728 1170
rect 5184 1142 5304 1170
rect 7760 1142 7880 1170
rect 2608 800 2636 1142
rect 5184 800 5212 1142
rect 7760 800 7788 1142
rect 10244 898 10272 2246
rect 10380 2204 10688 2213
rect 10380 2202 10386 2204
rect 10442 2202 10466 2204
rect 10522 2202 10546 2204
rect 10602 2202 10626 2204
rect 10682 2202 10688 2204
rect 10442 2150 10444 2202
rect 10624 2150 10626 2202
rect 10380 2148 10386 2150
rect 10442 2148 10466 2150
rect 10522 2148 10546 2150
rect 10602 2148 10626 2150
rect 10682 2148 10688 2150
rect 10380 2139 10688 2148
rect 13648 1306 13676 2382
rect 16224 1306 16252 2382
rect 18800 1306 18828 2382
rect 19810 2204 20118 2213
rect 19810 2202 19816 2204
rect 19872 2202 19896 2204
rect 19952 2202 19976 2204
rect 20032 2202 20056 2204
rect 20112 2202 20118 2204
rect 19872 2150 19874 2202
rect 20054 2150 20056 2202
rect 19810 2148 19816 2150
rect 19872 2148 19896 2150
rect 19952 2148 19976 2150
rect 20032 2148 20056 2150
rect 20112 2148 20118 2150
rect 19810 2139 20118 2148
rect 21376 1306 21404 2382
rect 23952 1306 23980 2382
rect 27172 1306 27200 2382
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 34888 2304 34940 2310
rect 34888 2246 34940 2252
rect 29240 2204 29548 2213
rect 29240 2202 29246 2204
rect 29302 2202 29326 2204
rect 29382 2202 29406 2204
rect 29462 2202 29486 2204
rect 29542 2202 29548 2204
rect 29302 2150 29304 2202
rect 29484 2150 29486 2202
rect 29240 2148 29246 2150
rect 29302 2148 29326 2150
rect 29382 2148 29406 2150
rect 29462 2148 29486 2150
rect 29542 2148 29548 2150
rect 29240 2139 29548 2148
rect 13556 1278 13676 1306
rect 16132 1278 16252 1306
rect 18708 1278 18828 1306
rect 21284 1278 21404 1306
rect 23860 1278 23980 1306
rect 27080 1278 27200 1306
rect 10244 870 10364 898
rect 10336 800 10364 870
rect 13556 800 13584 1278
rect 16132 800 16160 1278
rect 18708 800 18736 1278
rect 21284 800 21312 1278
rect 23860 800 23888 1278
rect 27080 800 27108 1278
rect 29748 1170 29776 2246
rect 32324 1170 32352 2246
rect 34900 1170 34928 2246
rect 37476 1306 37504 2382
rect 29656 1142 29776 1170
rect 32232 1142 32352 1170
rect 34808 1142 34928 1170
rect 37384 1278 37504 1306
rect 29656 800 29684 1142
rect 32232 800 32260 1142
rect 34808 800 34836 1142
rect 37384 800 37412 1278
rect 124 734 336 762
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 13542 0 13598 800
rect 16118 0 16174 800
rect 18694 0 18750 800
rect 21270 0 21326 800
rect 23846 0 23902 800
rect 27066 0 27122 800
rect 29642 0 29698 800
rect 32218 0 32274 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 38488 785 38516 2382
rect 38670 2204 38978 2213
rect 38670 2202 38676 2204
rect 38732 2202 38756 2204
rect 38812 2202 38836 2204
rect 38892 2202 38916 2204
rect 38972 2202 38978 2204
rect 38732 2150 38734 2202
rect 38914 2150 38916 2202
rect 38670 2148 38676 2150
rect 38732 2148 38756 2150
rect 38812 2148 38836 2150
rect 38892 2148 38916 2150
rect 38972 2148 38978 2150
rect 38670 2139 38978 2148
rect 38474 776 38530 785
rect 38474 711 38530 720
<< via2 >>
rect 2778 10920 2834 10976
rect 10386 9818 10442 9820
rect 10466 9818 10522 9820
rect 10546 9818 10602 9820
rect 10626 9818 10682 9820
rect 10386 9766 10432 9818
rect 10432 9766 10442 9818
rect 10466 9766 10496 9818
rect 10496 9766 10508 9818
rect 10508 9766 10522 9818
rect 10546 9766 10560 9818
rect 10560 9766 10572 9818
rect 10572 9766 10602 9818
rect 10626 9766 10636 9818
rect 10636 9766 10682 9818
rect 10386 9764 10442 9766
rect 10466 9764 10522 9766
rect 10546 9764 10602 9766
rect 10626 9764 10682 9766
rect 19816 9818 19872 9820
rect 19896 9818 19952 9820
rect 19976 9818 20032 9820
rect 20056 9818 20112 9820
rect 19816 9766 19862 9818
rect 19862 9766 19872 9818
rect 19896 9766 19926 9818
rect 19926 9766 19938 9818
rect 19938 9766 19952 9818
rect 19976 9766 19990 9818
rect 19990 9766 20002 9818
rect 20002 9766 20032 9818
rect 20056 9766 20066 9818
rect 20066 9766 20112 9818
rect 19816 9764 19872 9766
rect 19896 9764 19952 9766
rect 19976 9764 20032 9766
rect 20056 9764 20112 9766
rect 29246 9818 29302 9820
rect 29326 9818 29382 9820
rect 29406 9818 29462 9820
rect 29486 9818 29542 9820
rect 29246 9766 29292 9818
rect 29292 9766 29302 9818
rect 29326 9766 29356 9818
rect 29356 9766 29368 9818
rect 29368 9766 29382 9818
rect 29406 9766 29420 9818
rect 29420 9766 29432 9818
rect 29432 9766 29462 9818
rect 29486 9766 29496 9818
rect 29496 9766 29542 9818
rect 29246 9764 29302 9766
rect 29326 9764 29382 9766
rect 29406 9764 29462 9766
rect 29486 9764 29542 9766
rect 38676 9818 38732 9820
rect 38756 9818 38812 9820
rect 38836 9818 38892 9820
rect 38916 9818 38972 9820
rect 38676 9766 38722 9818
rect 38722 9766 38732 9818
rect 38756 9766 38786 9818
rect 38786 9766 38798 9818
rect 38798 9766 38812 9818
rect 38836 9766 38850 9818
rect 38850 9766 38862 9818
rect 38862 9766 38892 9818
rect 38916 9766 38926 9818
rect 38926 9766 38972 9818
rect 38676 9764 38732 9766
rect 38756 9764 38812 9766
rect 38836 9764 38892 9766
rect 38916 9764 38972 9766
rect 5671 9274 5727 9276
rect 5751 9274 5807 9276
rect 5831 9274 5887 9276
rect 5911 9274 5967 9276
rect 5671 9222 5717 9274
rect 5717 9222 5727 9274
rect 5751 9222 5781 9274
rect 5781 9222 5793 9274
rect 5793 9222 5807 9274
rect 5831 9222 5845 9274
rect 5845 9222 5857 9274
rect 5857 9222 5887 9274
rect 5911 9222 5921 9274
rect 5921 9222 5967 9274
rect 5671 9220 5727 9222
rect 5751 9220 5807 9222
rect 5831 9220 5887 9222
rect 5911 9220 5967 9222
rect 15101 9274 15157 9276
rect 15181 9274 15237 9276
rect 15261 9274 15317 9276
rect 15341 9274 15397 9276
rect 15101 9222 15147 9274
rect 15147 9222 15157 9274
rect 15181 9222 15211 9274
rect 15211 9222 15223 9274
rect 15223 9222 15237 9274
rect 15261 9222 15275 9274
rect 15275 9222 15287 9274
rect 15287 9222 15317 9274
rect 15341 9222 15351 9274
rect 15351 9222 15397 9274
rect 15101 9220 15157 9222
rect 15181 9220 15237 9222
rect 15261 9220 15317 9222
rect 15341 9220 15397 9222
rect 24531 9274 24587 9276
rect 24611 9274 24667 9276
rect 24691 9274 24747 9276
rect 24771 9274 24827 9276
rect 24531 9222 24577 9274
rect 24577 9222 24587 9274
rect 24611 9222 24641 9274
rect 24641 9222 24653 9274
rect 24653 9222 24667 9274
rect 24691 9222 24705 9274
rect 24705 9222 24717 9274
rect 24717 9222 24747 9274
rect 24771 9222 24781 9274
rect 24781 9222 24827 9274
rect 24531 9220 24587 9222
rect 24611 9220 24667 9222
rect 24691 9220 24747 9222
rect 24771 9220 24827 9222
rect 33961 9274 34017 9276
rect 34041 9274 34097 9276
rect 34121 9274 34177 9276
rect 34201 9274 34257 9276
rect 33961 9222 34007 9274
rect 34007 9222 34017 9274
rect 34041 9222 34071 9274
rect 34071 9222 34083 9274
rect 34083 9222 34097 9274
rect 34121 9222 34135 9274
rect 34135 9222 34147 9274
rect 34147 9222 34177 9274
rect 34201 9222 34211 9274
rect 34211 9222 34257 9274
rect 33961 9220 34017 9222
rect 34041 9220 34097 9222
rect 34121 9220 34177 9222
rect 34201 9220 34257 9222
rect 38474 8900 38530 8936
rect 38474 8880 38476 8900
rect 38476 8880 38528 8900
rect 38528 8880 38530 8900
rect 10386 8730 10442 8732
rect 10466 8730 10522 8732
rect 10546 8730 10602 8732
rect 10626 8730 10682 8732
rect 10386 8678 10432 8730
rect 10432 8678 10442 8730
rect 10466 8678 10496 8730
rect 10496 8678 10508 8730
rect 10508 8678 10522 8730
rect 10546 8678 10560 8730
rect 10560 8678 10572 8730
rect 10572 8678 10602 8730
rect 10626 8678 10636 8730
rect 10636 8678 10682 8730
rect 10386 8676 10442 8678
rect 10466 8676 10522 8678
rect 10546 8676 10602 8678
rect 10626 8676 10682 8678
rect 19816 8730 19872 8732
rect 19896 8730 19952 8732
rect 19976 8730 20032 8732
rect 20056 8730 20112 8732
rect 19816 8678 19862 8730
rect 19862 8678 19872 8730
rect 19896 8678 19926 8730
rect 19926 8678 19938 8730
rect 19938 8678 19952 8730
rect 19976 8678 19990 8730
rect 19990 8678 20002 8730
rect 20002 8678 20032 8730
rect 20056 8678 20066 8730
rect 20066 8678 20112 8730
rect 19816 8676 19872 8678
rect 19896 8676 19952 8678
rect 19976 8676 20032 8678
rect 20056 8676 20112 8678
rect 29246 8730 29302 8732
rect 29326 8730 29382 8732
rect 29406 8730 29462 8732
rect 29486 8730 29542 8732
rect 29246 8678 29292 8730
rect 29292 8678 29302 8730
rect 29326 8678 29356 8730
rect 29356 8678 29368 8730
rect 29368 8678 29382 8730
rect 29406 8678 29420 8730
rect 29420 8678 29432 8730
rect 29432 8678 29462 8730
rect 29486 8678 29496 8730
rect 29496 8678 29542 8730
rect 29246 8676 29302 8678
rect 29326 8676 29382 8678
rect 29406 8676 29462 8678
rect 29486 8676 29542 8678
rect 38676 8730 38732 8732
rect 38756 8730 38812 8732
rect 38836 8730 38892 8732
rect 38916 8730 38972 8732
rect 38676 8678 38722 8730
rect 38722 8678 38732 8730
rect 38756 8678 38786 8730
rect 38786 8678 38798 8730
rect 38798 8678 38812 8730
rect 38836 8678 38850 8730
rect 38850 8678 38862 8730
rect 38862 8678 38892 8730
rect 38916 8678 38926 8730
rect 38926 8678 38972 8730
rect 38676 8676 38732 8678
rect 38756 8676 38812 8678
rect 38836 8676 38892 8678
rect 38916 8676 38972 8678
rect 1398 8200 1454 8256
rect 5671 8186 5727 8188
rect 5751 8186 5807 8188
rect 5831 8186 5887 8188
rect 5911 8186 5967 8188
rect 5671 8134 5717 8186
rect 5717 8134 5727 8186
rect 5751 8134 5781 8186
rect 5781 8134 5793 8186
rect 5793 8134 5807 8186
rect 5831 8134 5845 8186
rect 5845 8134 5857 8186
rect 5857 8134 5887 8186
rect 5911 8134 5921 8186
rect 5921 8134 5967 8186
rect 5671 8132 5727 8134
rect 5751 8132 5807 8134
rect 5831 8132 5887 8134
rect 5911 8132 5967 8134
rect 15101 8186 15157 8188
rect 15181 8186 15237 8188
rect 15261 8186 15317 8188
rect 15341 8186 15397 8188
rect 15101 8134 15147 8186
rect 15147 8134 15157 8186
rect 15181 8134 15211 8186
rect 15211 8134 15223 8186
rect 15223 8134 15237 8186
rect 15261 8134 15275 8186
rect 15275 8134 15287 8186
rect 15287 8134 15317 8186
rect 15341 8134 15351 8186
rect 15351 8134 15397 8186
rect 15101 8132 15157 8134
rect 15181 8132 15237 8134
rect 15261 8132 15317 8134
rect 15341 8132 15397 8134
rect 24531 8186 24587 8188
rect 24611 8186 24667 8188
rect 24691 8186 24747 8188
rect 24771 8186 24827 8188
rect 24531 8134 24577 8186
rect 24577 8134 24587 8186
rect 24611 8134 24641 8186
rect 24641 8134 24653 8186
rect 24653 8134 24667 8186
rect 24691 8134 24705 8186
rect 24705 8134 24717 8186
rect 24717 8134 24747 8186
rect 24771 8134 24781 8186
rect 24781 8134 24827 8186
rect 24531 8132 24587 8134
rect 24611 8132 24667 8134
rect 24691 8132 24747 8134
rect 24771 8132 24827 8134
rect 33961 8186 34017 8188
rect 34041 8186 34097 8188
rect 34121 8186 34177 8188
rect 34201 8186 34257 8188
rect 33961 8134 34007 8186
rect 34007 8134 34017 8186
rect 34041 8134 34071 8186
rect 34071 8134 34083 8186
rect 34083 8134 34097 8186
rect 34121 8134 34135 8186
rect 34135 8134 34147 8186
rect 34147 8134 34177 8186
rect 34201 8134 34211 8186
rect 34211 8134 34257 8186
rect 33961 8132 34017 8134
rect 34041 8132 34097 8134
rect 34121 8132 34177 8134
rect 34201 8132 34257 8134
rect 10386 7642 10442 7644
rect 10466 7642 10522 7644
rect 10546 7642 10602 7644
rect 10626 7642 10682 7644
rect 10386 7590 10432 7642
rect 10432 7590 10442 7642
rect 10466 7590 10496 7642
rect 10496 7590 10508 7642
rect 10508 7590 10522 7642
rect 10546 7590 10560 7642
rect 10560 7590 10572 7642
rect 10572 7590 10602 7642
rect 10626 7590 10636 7642
rect 10636 7590 10682 7642
rect 10386 7588 10442 7590
rect 10466 7588 10522 7590
rect 10546 7588 10602 7590
rect 10626 7588 10682 7590
rect 19816 7642 19872 7644
rect 19896 7642 19952 7644
rect 19976 7642 20032 7644
rect 20056 7642 20112 7644
rect 19816 7590 19862 7642
rect 19862 7590 19872 7642
rect 19896 7590 19926 7642
rect 19926 7590 19938 7642
rect 19938 7590 19952 7642
rect 19976 7590 19990 7642
rect 19990 7590 20002 7642
rect 20002 7590 20032 7642
rect 20056 7590 20066 7642
rect 20066 7590 20112 7642
rect 19816 7588 19872 7590
rect 19896 7588 19952 7590
rect 19976 7588 20032 7590
rect 20056 7588 20112 7590
rect 29246 7642 29302 7644
rect 29326 7642 29382 7644
rect 29406 7642 29462 7644
rect 29486 7642 29542 7644
rect 29246 7590 29292 7642
rect 29292 7590 29302 7642
rect 29326 7590 29356 7642
rect 29356 7590 29368 7642
rect 29368 7590 29382 7642
rect 29406 7590 29420 7642
rect 29420 7590 29432 7642
rect 29432 7590 29462 7642
rect 29486 7590 29496 7642
rect 29496 7590 29542 7642
rect 29246 7588 29302 7590
rect 29326 7588 29382 7590
rect 29406 7588 29462 7590
rect 29486 7588 29542 7590
rect 38676 7642 38732 7644
rect 38756 7642 38812 7644
rect 38836 7642 38892 7644
rect 38916 7642 38972 7644
rect 38676 7590 38722 7642
rect 38722 7590 38732 7642
rect 38756 7590 38786 7642
rect 38786 7590 38798 7642
rect 38798 7590 38812 7642
rect 38836 7590 38850 7642
rect 38850 7590 38862 7642
rect 38862 7590 38892 7642
rect 38916 7590 38926 7642
rect 38926 7590 38972 7642
rect 38676 7588 38732 7590
rect 38756 7588 38812 7590
rect 38836 7588 38892 7590
rect 38916 7588 38972 7590
rect 5671 7098 5727 7100
rect 5751 7098 5807 7100
rect 5831 7098 5887 7100
rect 5911 7098 5967 7100
rect 5671 7046 5717 7098
rect 5717 7046 5727 7098
rect 5751 7046 5781 7098
rect 5781 7046 5793 7098
rect 5793 7046 5807 7098
rect 5831 7046 5845 7098
rect 5845 7046 5857 7098
rect 5857 7046 5887 7098
rect 5911 7046 5921 7098
rect 5921 7046 5967 7098
rect 5671 7044 5727 7046
rect 5751 7044 5807 7046
rect 5831 7044 5887 7046
rect 5911 7044 5967 7046
rect 15101 7098 15157 7100
rect 15181 7098 15237 7100
rect 15261 7098 15317 7100
rect 15341 7098 15397 7100
rect 15101 7046 15147 7098
rect 15147 7046 15157 7098
rect 15181 7046 15211 7098
rect 15211 7046 15223 7098
rect 15223 7046 15237 7098
rect 15261 7046 15275 7098
rect 15275 7046 15287 7098
rect 15287 7046 15317 7098
rect 15341 7046 15351 7098
rect 15351 7046 15397 7098
rect 15101 7044 15157 7046
rect 15181 7044 15237 7046
rect 15261 7044 15317 7046
rect 15341 7044 15397 7046
rect 24531 7098 24587 7100
rect 24611 7098 24667 7100
rect 24691 7098 24747 7100
rect 24771 7098 24827 7100
rect 24531 7046 24577 7098
rect 24577 7046 24587 7098
rect 24611 7046 24641 7098
rect 24641 7046 24653 7098
rect 24653 7046 24667 7098
rect 24691 7046 24705 7098
rect 24705 7046 24717 7098
rect 24717 7046 24747 7098
rect 24771 7046 24781 7098
rect 24781 7046 24827 7098
rect 24531 7044 24587 7046
rect 24611 7044 24667 7046
rect 24691 7044 24747 7046
rect 24771 7044 24827 7046
rect 33961 7098 34017 7100
rect 34041 7098 34097 7100
rect 34121 7098 34177 7100
rect 34201 7098 34257 7100
rect 33961 7046 34007 7098
rect 34007 7046 34017 7098
rect 34041 7046 34071 7098
rect 34071 7046 34083 7098
rect 34083 7046 34097 7098
rect 34121 7046 34135 7098
rect 34135 7046 34147 7098
rect 34147 7046 34177 7098
rect 34201 7046 34211 7098
rect 34211 7046 34257 7098
rect 33961 7044 34017 7046
rect 34041 7044 34097 7046
rect 34121 7044 34177 7046
rect 34201 7044 34257 7046
rect 10386 6554 10442 6556
rect 10466 6554 10522 6556
rect 10546 6554 10602 6556
rect 10626 6554 10682 6556
rect 10386 6502 10432 6554
rect 10432 6502 10442 6554
rect 10466 6502 10496 6554
rect 10496 6502 10508 6554
rect 10508 6502 10522 6554
rect 10546 6502 10560 6554
rect 10560 6502 10572 6554
rect 10572 6502 10602 6554
rect 10626 6502 10636 6554
rect 10636 6502 10682 6554
rect 10386 6500 10442 6502
rect 10466 6500 10522 6502
rect 10546 6500 10602 6502
rect 10626 6500 10682 6502
rect 19816 6554 19872 6556
rect 19896 6554 19952 6556
rect 19976 6554 20032 6556
rect 20056 6554 20112 6556
rect 19816 6502 19862 6554
rect 19862 6502 19872 6554
rect 19896 6502 19926 6554
rect 19926 6502 19938 6554
rect 19938 6502 19952 6554
rect 19976 6502 19990 6554
rect 19990 6502 20002 6554
rect 20002 6502 20032 6554
rect 20056 6502 20066 6554
rect 20066 6502 20112 6554
rect 19816 6500 19872 6502
rect 19896 6500 19952 6502
rect 19976 6500 20032 6502
rect 20056 6500 20112 6502
rect 29246 6554 29302 6556
rect 29326 6554 29382 6556
rect 29406 6554 29462 6556
rect 29486 6554 29542 6556
rect 29246 6502 29292 6554
rect 29292 6502 29302 6554
rect 29326 6502 29356 6554
rect 29356 6502 29368 6554
rect 29368 6502 29382 6554
rect 29406 6502 29420 6554
rect 29420 6502 29432 6554
rect 29432 6502 29462 6554
rect 29486 6502 29496 6554
rect 29496 6502 29542 6554
rect 29246 6500 29302 6502
rect 29326 6500 29382 6502
rect 29406 6500 29462 6502
rect 29486 6500 29542 6502
rect 38676 6554 38732 6556
rect 38756 6554 38812 6556
rect 38836 6554 38892 6556
rect 38916 6554 38972 6556
rect 38676 6502 38722 6554
rect 38722 6502 38732 6554
rect 38756 6502 38786 6554
rect 38786 6502 38798 6554
rect 38798 6502 38812 6554
rect 38836 6502 38850 6554
rect 38850 6502 38862 6554
rect 38862 6502 38892 6554
rect 38916 6502 38926 6554
rect 38926 6502 38972 6554
rect 38676 6500 38732 6502
rect 38756 6500 38812 6502
rect 38836 6500 38892 6502
rect 38916 6500 38972 6502
rect 38474 6196 38476 6216
rect 38476 6196 38528 6216
rect 38528 6196 38530 6216
rect 38474 6160 38530 6196
rect 5671 6010 5727 6012
rect 5751 6010 5807 6012
rect 5831 6010 5887 6012
rect 5911 6010 5967 6012
rect 5671 5958 5717 6010
rect 5717 5958 5727 6010
rect 5751 5958 5781 6010
rect 5781 5958 5793 6010
rect 5793 5958 5807 6010
rect 5831 5958 5845 6010
rect 5845 5958 5857 6010
rect 5857 5958 5887 6010
rect 5911 5958 5921 6010
rect 5921 5958 5967 6010
rect 5671 5956 5727 5958
rect 5751 5956 5807 5958
rect 5831 5956 5887 5958
rect 5911 5956 5967 5958
rect 15101 6010 15157 6012
rect 15181 6010 15237 6012
rect 15261 6010 15317 6012
rect 15341 6010 15397 6012
rect 15101 5958 15147 6010
rect 15147 5958 15157 6010
rect 15181 5958 15211 6010
rect 15211 5958 15223 6010
rect 15223 5958 15237 6010
rect 15261 5958 15275 6010
rect 15275 5958 15287 6010
rect 15287 5958 15317 6010
rect 15341 5958 15351 6010
rect 15351 5958 15397 6010
rect 15101 5956 15157 5958
rect 15181 5956 15237 5958
rect 15261 5956 15317 5958
rect 15341 5956 15397 5958
rect 24531 6010 24587 6012
rect 24611 6010 24667 6012
rect 24691 6010 24747 6012
rect 24771 6010 24827 6012
rect 24531 5958 24577 6010
rect 24577 5958 24587 6010
rect 24611 5958 24641 6010
rect 24641 5958 24653 6010
rect 24653 5958 24667 6010
rect 24691 5958 24705 6010
rect 24705 5958 24717 6010
rect 24717 5958 24747 6010
rect 24771 5958 24781 6010
rect 24781 5958 24827 6010
rect 24531 5956 24587 5958
rect 24611 5956 24667 5958
rect 24691 5956 24747 5958
rect 24771 5956 24827 5958
rect 33961 6010 34017 6012
rect 34041 6010 34097 6012
rect 34121 6010 34177 6012
rect 34201 6010 34257 6012
rect 33961 5958 34007 6010
rect 34007 5958 34017 6010
rect 34041 5958 34071 6010
rect 34071 5958 34083 6010
rect 34083 5958 34097 6010
rect 34121 5958 34135 6010
rect 34135 5958 34147 6010
rect 34147 5958 34177 6010
rect 34201 5958 34211 6010
rect 34211 5958 34257 6010
rect 33961 5956 34017 5958
rect 34041 5956 34097 5958
rect 34121 5956 34177 5958
rect 34201 5956 34257 5958
rect 1398 5516 1400 5536
rect 1400 5516 1452 5536
rect 1452 5516 1454 5536
rect 1398 5480 1454 5516
rect 10386 5466 10442 5468
rect 10466 5466 10522 5468
rect 10546 5466 10602 5468
rect 10626 5466 10682 5468
rect 10386 5414 10432 5466
rect 10432 5414 10442 5466
rect 10466 5414 10496 5466
rect 10496 5414 10508 5466
rect 10508 5414 10522 5466
rect 10546 5414 10560 5466
rect 10560 5414 10572 5466
rect 10572 5414 10602 5466
rect 10626 5414 10636 5466
rect 10636 5414 10682 5466
rect 10386 5412 10442 5414
rect 10466 5412 10522 5414
rect 10546 5412 10602 5414
rect 10626 5412 10682 5414
rect 19816 5466 19872 5468
rect 19896 5466 19952 5468
rect 19976 5466 20032 5468
rect 20056 5466 20112 5468
rect 19816 5414 19862 5466
rect 19862 5414 19872 5466
rect 19896 5414 19926 5466
rect 19926 5414 19938 5466
rect 19938 5414 19952 5466
rect 19976 5414 19990 5466
rect 19990 5414 20002 5466
rect 20002 5414 20032 5466
rect 20056 5414 20066 5466
rect 20066 5414 20112 5466
rect 19816 5412 19872 5414
rect 19896 5412 19952 5414
rect 19976 5412 20032 5414
rect 20056 5412 20112 5414
rect 29246 5466 29302 5468
rect 29326 5466 29382 5468
rect 29406 5466 29462 5468
rect 29486 5466 29542 5468
rect 29246 5414 29292 5466
rect 29292 5414 29302 5466
rect 29326 5414 29356 5466
rect 29356 5414 29368 5466
rect 29368 5414 29382 5466
rect 29406 5414 29420 5466
rect 29420 5414 29432 5466
rect 29432 5414 29462 5466
rect 29486 5414 29496 5466
rect 29496 5414 29542 5466
rect 29246 5412 29302 5414
rect 29326 5412 29382 5414
rect 29406 5412 29462 5414
rect 29486 5412 29542 5414
rect 38676 5466 38732 5468
rect 38756 5466 38812 5468
rect 38836 5466 38892 5468
rect 38916 5466 38972 5468
rect 38676 5414 38722 5466
rect 38722 5414 38732 5466
rect 38756 5414 38786 5466
rect 38786 5414 38798 5466
rect 38798 5414 38812 5466
rect 38836 5414 38850 5466
rect 38850 5414 38862 5466
rect 38862 5414 38892 5466
rect 38916 5414 38926 5466
rect 38926 5414 38972 5466
rect 38676 5412 38732 5414
rect 38756 5412 38812 5414
rect 38836 5412 38892 5414
rect 38916 5412 38972 5414
rect 5671 4922 5727 4924
rect 5751 4922 5807 4924
rect 5831 4922 5887 4924
rect 5911 4922 5967 4924
rect 5671 4870 5717 4922
rect 5717 4870 5727 4922
rect 5751 4870 5781 4922
rect 5781 4870 5793 4922
rect 5793 4870 5807 4922
rect 5831 4870 5845 4922
rect 5845 4870 5857 4922
rect 5857 4870 5887 4922
rect 5911 4870 5921 4922
rect 5921 4870 5967 4922
rect 5671 4868 5727 4870
rect 5751 4868 5807 4870
rect 5831 4868 5887 4870
rect 5911 4868 5967 4870
rect 15101 4922 15157 4924
rect 15181 4922 15237 4924
rect 15261 4922 15317 4924
rect 15341 4922 15397 4924
rect 15101 4870 15147 4922
rect 15147 4870 15157 4922
rect 15181 4870 15211 4922
rect 15211 4870 15223 4922
rect 15223 4870 15237 4922
rect 15261 4870 15275 4922
rect 15275 4870 15287 4922
rect 15287 4870 15317 4922
rect 15341 4870 15351 4922
rect 15351 4870 15397 4922
rect 15101 4868 15157 4870
rect 15181 4868 15237 4870
rect 15261 4868 15317 4870
rect 15341 4868 15397 4870
rect 24531 4922 24587 4924
rect 24611 4922 24667 4924
rect 24691 4922 24747 4924
rect 24771 4922 24827 4924
rect 24531 4870 24577 4922
rect 24577 4870 24587 4922
rect 24611 4870 24641 4922
rect 24641 4870 24653 4922
rect 24653 4870 24667 4922
rect 24691 4870 24705 4922
rect 24705 4870 24717 4922
rect 24717 4870 24747 4922
rect 24771 4870 24781 4922
rect 24781 4870 24827 4922
rect 24531 4868 24587 4870
rect 24611 4868 24667 4870
rect 24691 4868 24747 4870
rect 24771 4868 24827 4870
rect 33961 4922 34017 4924
rect 34041 4922 34097 4924
rect 34121 4922 34177 4924
rect 34201 4922 34257 4924
rect 33961 4870 34007 4922
rect 34007 4870 34017 4922
rect 34041 4870 34071 4922
rect 34071 4870 34083 4922
rect 34083 4870 34097 4922
rect 34121 4870 34135 4922
rect 34135 4870 34147 4922
rect 34147 4870 34177 4922
rect 34201 4870 34211 4922
rect 34211 4870 34257 4922
rect 33961 4868 34017 4870
rect 34041 4868 34097 4870
rect 34121 4868 34177 4870
rect 34201 4868 34257 4870
rect 10386 4378 10442 4380
rect 10466 4378 10522 4380
rect 10546 4378 10602 4380
rect 10626 4378 10682 4380
rect 10386 4326 10432 4378
rect 10432 4326 10442 4378
rect 10466 4326 10496 4378
rect 10496 4326 10508 4378
rect 10508 4326 10522 4378
rect 10546 4326 10560 4378
rect 10560 4326 10572 4378
rect 10572 4326 10602 4378
rect 10626 4326 10636 4378
rect 10636 4326 10682 4378
rect 10386 4324 10442 4326
rect 10466 4324 10522 4326
rect 10546 4324 10602 4326
rect 10626 4324 10682 4326
rect 19816 4378 19872 4380
rect 19896 4378 19952 4380
rect 19976 4378 20032 4380
rect 20056 4378 20112 4380
rect 19816 4326 19862 4378
rect 19862 4326 19872 4378
rect 19896 4326 19926 4378
rect 19926 4326 19938 4378
rect 19938 4326 19952 4378
rect 19976 4326 19990 4378
rect 19990 4326 20002 4378
rect 20002 4326 20032 4378
rect 20056 4326 20066 4378
rect 20066 4326 20112 4378
rect 19816 4324 19872 4326
rect 19896 4324 19952 4326
rect 19976 4324 20032 4326
rect 20056 4324 20112 4326
rect 29246 4378 29302 4380
rect 29326 4378 29382 4380
rect 29406 4378 29462 4380
rect 29486 4378 29542 4380
rect 29246 4326 29292 4378
rect 29292 4326 29302 4378
rect 29326 4326 29356 4378
rect 29356 4326 29368 4378
rect 29368 4326 29382 4378
rect 29406 4326 29420 4378
rect 29420 4326 29432 4378
rect 29432 4326 29462 4378
rect 29486 4326 29496 4378
rect 29496 4326 29542 4378
rect 29246 4324 29302 4326
rect 29326 4324 29382 4326
rect 29406 4324 29462 4326
rect 29486 4324 29542 4326
rect 38676 4378 38732 4380
rect 38756 4378 38812 4380
rect 38836 4378 38892 4380
rect 38916 4378 38972 4380
rect 38676 4326 38722 4378
rect 38722 4326 38732 4378
rect 38756 4326 38786 4378
rect 38786 4326 38798 4378
rect 38798 4326 38812 4378
rect 38836 4326 38850 4378
rect 38850 4326 38862 4378
rect 38862 4326 38892 4378
rect 38916 4326 38926 4378
rect 38926 4326 38972 4378
rect 38676 4324 38732 4326
rect 38756 4324 38812 4326
rect 38836 4324 38892 4326
rect 38916 4324 38972 4326
rect 5671 3834 5727 3836
rect 5751 3834 5807 3836
rect 5831 3834 5887 3836
rect 5911 3834 5967 3836
rect 5671 3782 5717 3834
rect 5717 3782 5727 3834
rect 5751 3782 5781 3834
rect 5781 3782 5793 3834
rect 5793 3782 5807 3834
rect 5831 3782 5845 3834
rect 5845 3782 5857 3834
rect 5857 3782 5887 3834
rect 5911 3782 5921 3834
rect 5921 3782 5967 3834
rect 5671 3780 5727 3782
rect 5751 3780 5807 3782
rect 5831 3780 5887 3782
rect 5911 3780 5967 3782
rect 15101 3834 15157 3836
rect 15181 3834 15237 3836
rect 15261 3834 15317 3836
rect 15341 3834 15397 3836
rect 15101 3782 15147 3834
rect 15147 3782 15157 3834
rect 15181 3782 15211 3834
rect 15211 3782 15223 3834
rect 15223 3782 15237 3834
rect 15261 3782 15275 3834
rect 15275 3782 15287 3834
rect 15287 3782 15317 3834
rect 15341 3782 15351 3834
rect 15351 3782 15397 3834
rect 15101 3780 15157 3782
rect 15181 3780 15237 3782
rect 15261 3780 15317 3782
rect 15341 3780 15397 3782
rect 24531 3834 24587 3836
rect 24611 3834 24667 3836
rect 24691 3834 24747 3836
rect 24771 3834 24827 3836
rect 24531 3782 24577 3834
rect 24577 3782 24587 3834
rect 24611 3782 24641 3834
rect 24641 3782 24653 3834
rect 24653 3782 24667 3834
rect 24691 3782 24705 3834
rect 24705 3782 24717 3834
rect 24717 3782 24747 3834
rect 24771 3782 24781 3834
rect 24781 3782 24827 3834
rect 24531 3780 24587 3782
rect 24611 3780 24667 3782
rect 24691 3780 24747 3782
rect 24771 3780 24827 3782
rect 33961 3834 34017 3836
rect 34041 3834 34097 3836
rect 34121 3834 34177 3836
rect 34201 3834 34257 3836
rect 33961 3782 34007 3834
rect 34007 3782 34017 3834
rect 34041 3782 34071 3834
rect 34071 3782 34083 3834
rect 34083 3782 34097 3834
rect 34121 3782 34135 3834
rect 34135 3782 34147 3834
rect 34147 3782 34177 3834
rect 34201 3782 34211 3834
rect 34211 3782 34257 3834
rect 33961 3780 34017 3782
rect 34041 3780 34097 3782
rect 34121 3780 34177 3782
rect 34201 3780 34257 3782
rect 38474 3476 38476 3496
rect 38476 3476 38528 3496
rect 38528 3476 38530 3496
rect 38474 3440 38530 3476
rect 10386 3290 10442 3292
rect 10466 3290 10522 3292
rect 10546 3290 10602 3292
rect 10626 3290 10682 3292
rect 10386 3238 10432 3290
rect 10432 3238 10442 3290
rect 10466 3238 10496 3290
rect 10496 3238 10508 3290
rect 10508 3238 10522 3290
rect 10546 3238 10560 3290
rect 10560 3238 10572 3290
rect 10572 3238 10602 3290
rect 10626 3238 10636 3290
rect 10636 3238 10682 3290
rect 10386 3236 10442 3238
rect 10466 3236 10522 3238
rect 10546 3236 10602 3238
rect 10626 3236 10682 3238
rect 19816 3290 19872 3292
rect 19896 3290 19952 3292
rect 19976 3290 20032 3292
rect 20056 3290 20112 3292
rect 19816 3238 19862 3290
rect 19862 3238 19872 3290
rect 19896 3238 19926 3290
rect 19926 3238 19938 3290
rect 19938 3238 19952 3290
rect 19976 3238 19990 3290
rect 19990 3238 20002 3290
rect 20002 3238 20032 3290
rect 20056 3238 20066 3290
rect 20066 3238 20112 3290
rect 19816 3236 19872 3238
rect 19896 3236 19952 3238
rect 19976 3236 20032 3238
rect 20056 3236 20112 3238
rect 29246 3290 29302 3292
rect 29326 3290 29382 3292
rect 29406 3290 29462 3292
rect 29486 3290 29542 3292
rect 29246 3238 29292 3290
rect 29292 3238 29302 3290
rect 29326 3238 29356 3290
rect 29356 3238 29368 3290
rect 29368 3238 29382 3290
rect 29406 3238 29420 3290
rect 29420 3238 29432 3290
rect 29432 3238 29462 3290
rect 29486 3238 29496 3290
rect 29496 3238 29542 3290
rect 29246 3236 29302 3238
rect 29326 3236 29382 3238
rect 29406 3236 29462 3238
rect 29486 3236 29542 3238
rect 38676 3290 38732 3292
rect 38756 3290 38812 3292
rect 38836 3290 38892 3292
rect 38916 3290 38972 3292
rect 38676 3238 38722 3290
rect 38722 3238 38732 3290
rect 38756 3238 38786 3290
rect 38786 3238 38798 3290
rect 38798 3238 38812 3290
rect 38836 3238 38850 3290
rect 38850 3238 38862 3290
rect 38862 3238 38892 3290
rect 38916 3238 38926 3290
rect 38926 3238 38972 3290
rect 38676 3236 38732 3238
rect 38756 3236 38812 3238
rect 38836 3236 38892 3238
rect 38916 3236 38972 3238
rect 938 2760 994 2816
rect 5671 2746 5727 2748
rect 5751 2746 5807 2748
rect 5831 2746 5887 2748
rect 5911 2746 5967 2748
rect 5671 2694 5717 2746
rect 5717 2694 5727 2746
rect 5751 2694 5781 2746
rect 5781 2694 5793 2746
rect 5793 2694 5807 2746
rect 5831 2694 5845 2746
rect 5845 2694 5857 2746
rect 5857 2694 5887 2746
rect 5911 2694 5921 2746
rect 5921 2694 5967 2746
rect 5671 2692 5727 2694
rect 5751 2692 5807 2694
rect 5831 2692 5887 2694
rect 5911 2692 5967 2694
rect 15101 2746 15157 2748
rect 15181 2746 15237 2748
rect 15261 2746 15317 2748
rect 15341 2746 15397 2748
rect 15101 2694 15147 2746
rect 15147 2694 15157 2746
rect 15181 2694 15211 2746
rect 15211 2694 15223 2746
rect 15223 2694 15237 2746
rect 15261 2694 15275 2746
rect 15275 2694 15287 2746
rect 15287 2694 15317 2746
rect 15341 2694 15351 2746
rect 15351 2694 15397 2746
rect 15101 2692 15157 2694
rect 15181 2692 15237 2694
rect 15261 2692 15317 2694
rect 15341 2692 15397 2694
rect 24531 2746 24587 2748
rect 24611 2746 24667 2748
rect 24691 2746 24747 2748
rect 24771 2746 24827 2748
rect 24531 2694 24577 2746
rect 24577 2694 24587 2746
rect 24611 2694 24641 2746
rect 24641 2694 24653 2746
rect 24653 2694 24667 2746
rect 24691 2694 24705 2746
rect 24705 2694 24717 2746
rect 24717 2694 24747 2746
rect 24771 2694 24781 2746
rect 24781 2694 24827 2746
rect 24531 2692 24587 2694
rect 24611 2692 24667 2694
rect 24691 2692 24747 2694
rect 24771 2692 24827 2694
rect 33961 2746 34017 2748
rect 34041 2746 34097 2748
rect 34121 2746 34177 2748
rect 34201 2746 34257 2748
rect 33961 2694 34007 2746
rect 34007 2694 34017 2746
rect 34041 2694 34071 2746
rect 34071 2694 34083 2746
rect 34083 2694 34097 2746
rect 34121 2694 34135 2746
rect 34135 2694 34147 2746
rect 34147 2694 34177 2746
rect 34201 2694 34211 2746
rect 34211 2694 34257 2746
rect 33961 2692 34017 2694
rect 34041 2692 34097 2694
rect 34121 2692 34177 2694
rect 34201 2692 34257 2694
rect 10386 2202 10442 2204
rect 10466 2202 10522 2204
rect 10546 2202 10602 2204
rect 10626 2202 10682 2204
rect 10386 2150 10432 2202
rect 10432 2150 10442 2202
rect 10466 2150 10496 2202
rect 10496 2150 10508 2202
rect 10508 2150 10522 2202
rect 10546 2150 10560 2202
rect 10560 2150 10572 2202
rect 10572 2150 10602 2202
rect 10626 2150 10636 2202
rect 10636 2150 10682 2202
rect 10386 2148 10442 2150
rect 10466 2148 10522 2150
rect 10546 2148 10602 2150
rect 10626 2148 10682 2150
rect 19816 2202 19872 2204
rect 19896 2202 19952 2204
rect 19976 2202 20032 2204
rect 20056 2202 20112 2204
rect 19816 2150 19862 2202
rect 19862 2150 19872 2202
rect 19896 2150 19926 2202
rect 19926 2150 19938 2202
rect 19938 2150 19952 2202
rect 19976 2150 19990 2202
rect 19990 2150 20002 2202
rect 20002 2150 20032 2202
rect 20056 2150 20066 2202
rect 20066 2150 20112 2202
rect 19816 2148 19872 2150
rect 19896 2148 19952 2150
rect 19976 2148 20032 2150
rect 20056 2148 20112 2150
rect 29246 2202 29302 2204
rect 29326 2202 29382 2204
rect 29406 2202 29462 2204
rect 29486 2202 29542 2204
rect 29246 2150 29292 2202
rect 29292 2150 29302 2202
rect 29326 2150 29356 2202
rect 29356 2150 29368 2202
rect 29368 2150 29382 2202
rect 29406 2150 29420 2202
rect 29420 2150 29432 2202
rect 29432 2150 29462 2202
rect 29486 2150 29496 2202
rect 29496 2150 29542 2202
rect 29246 2148 29302 2150
rect 29326 2148 29382 2150
rect 29406 2148 29462 2150
rect 29486 2148 29542 2150
rect 38676 2202 38732 2204
rect 38756 2202 38812 2204
rect 38836 2202 38892 2204
rect 38916 2202 38972 2204
rect 38676 2150 38722 2202
rect 38722 2150 38732 2202
rect 38756 2150 38786 2202
rect 38786 2150 38798 2202
rect 38798 2150 38812 2202
rect 38836 2150 38850 2202
rect 38850 2150 38862 2202
rect 38862 2150 38892 2202
rect 38916 2150 38926 2202
rect 38926 2150 38972 2202
rect 38676 2148 38732 2150
rect 38756 2148 38812 2150
rect 38836 2148 38892 2150
rect 38916 2148 38972 2150
rect 38474 720 38530 776
<< metal3 >>
rect 0 10978 800 11008
rect 2773 10978 2839 10981
rect 0 10976 2839 10978
rect 0 10920 2778 10976
rect 2834 10920 2839 10976
rect 0 10918 2839 10920
rect 0 10888 800 10918
rect 2773 10915 2839 10918
rect 10376 9824 10692 9825
rect 10376 9760 10382 9824
rect 10446 9760 10462 9824
rect 10526 9760 10542 9824
rect 10606 9760 10622 9824
rect 10686 9760 10692 9824
rect 10376 9759 10692 9760
rect 19806 9824 20122 9825
rect 19806 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20052 9824
rect 20116 9760 20122 9824
rect 19806 9759 20122 9760
rect 29236 9824 29552 9825
rect 29236 9760 29242 9824
rect 29306 9760 29322 9824
rect 29386 9760 29402 9824
rect 29466 9760 29482 9824
rect 29546 9760 29552 9824
rect 29236 9759 29552 9760
rect 38666 9824 38982 9825
rect 38666 9760 38672 9824
rect 38736 9760 38752 9824
rect 38816 9760 38832 9824
rect 38896 9760 38912 9824
rect 38976 9760 38982 9824
rect 38666 9759 38982 9760
rect 5661 9280 5977 9281
rect 5661 9216 5667 9280
rect 5731 9216 5747 9280
rect 5811 9216 5827 9280
rect 5891 9216 5907 9280
rect 5971 9216 5977 9280
rect 5661 9215 5977 9216
rect 15091 9280 15407 9281
rect 15091 9216 15097 9280
rect 15161 9216 15177 9280
rect 15241 9216 15257 9280
rect 15321 9216 15337 9280
rect 15401 9216 15407 9280
rect 15091 9215 15407 9216
rect 24521 9280 24837 9281
rect 24521 9216 24527 9280
rect 24591 9216 24607 9280
rect 24671 9216 24687 9280
rect 24751 9216 24767 9280
rect 24831 9216 24837 9280
rect 24521 9215 24837 9216
rect 33951 9280 34267 9281
rect 33951 9216 33957 9280
rect 34021 9216 34037 9280
rect 34101 9216 34117 9280
rect 34181 9216 34197 9280
rect 34261 9216 34267 9280
rect 33951 9215 34267 9216
rect 38469 8938 38535 8941
rect 39200 8938 40000 8968
rect 38469 8936 40000 8938
rect 38469 8880 38474 8936
rect 38530 8880 40000 8936
rect 38469 8878 40000 8880
rect 38469 8875 38535 8878
rect 39200 8848 40000 8878
rect 10376 8736 10692 8737
rect 10376 8672 10382 8736
rect 10446 8672 10462 8736
rect 10526 8672 10542 8736
rect 10606 8672 10622 8736
rect 10686 8672 10692 8736
rect 10376 8671 10692 8672
rect 19806 8736 20122 8737
rect 19806 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20052 8736
rect 20116 8672 20122 8736
rect 19806 8671 20122 8672
rect 29236 8736 29552 8737
rect 29236 8672 29242 8736
rect 29306 8672 29322 8736
rect 29386 8672 29402 8736
rect 29466 8672 29482 8736
rect 29546 8672 29552 8736
rect 29236 8671 29552 8672
rect 38666 8736 38982 8737
rect 38666 8672 38672 8736
rect 38736 8672 38752 8736
rect 38816 8672 38832 8736
rect 38896 8672 38912 8736
rect 38976 8672 38982 8736
rect 38666 8671 38982 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 5661 8192 5977 8193
rect 5661 8128 5667 8192
rect 5731 8128 5747 8192
rect 5811 8128 5827 8192
rect 5891 8128 5907 8192
rect 5971 8128 5977 8192
rect 5661 8127 5977 8128
rect 15091 8192 15407 8193
rect 15091 8128 15097 8192
rect 15161 8128 15177 8192
rect 15241 8128 15257 8192
rect 15321 8128 15337 8192
rect 15401 8128 15407 8192
rect 15091 8127 15407 8128
rect 24521 8192 24837 8193
rect 24521 8128 24527 8192
rect 24591 8128 24607 8192
rect 24671 8128 24687 8192
rect 24751 8128 24767 8192
rect 24831 8128 24837 8192
rect 24521 8127 24837 8128
rect 33951 8192 34267 8193
rect 33951 8128 33957 8192
rect 34021 8128 34037 8192
rect 34101 8128 34117 8192
rect 34181 8128 34197 8192
rect 34261 8128 34267 8192
rect 33951 8127 34267 8128
rect 10376 7648 10692 7649
rect 10376 7584 10382 7648
rect 10446 7584 10462 7648
rect 10526 7584 10542 7648
rect 10606 7584 10622 7648
rect 10686 7584 10692 7648
rect 10376 7583 10692 7584
rect 19806 7648 20122 7649
rect 19806 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20052 7648
rect 20116 7584 20122 7648
rect 19806 7583 20122 7584
rect 29236 7648 29552 7649
rect 29236 7584 29242 7648
rect 29306 7584 29322 7648
rect 29386 7584 29402 7648
rect 29466 7584 29482 7648
rect 29546 7584 29552 7648
rect 29236 7583 29552 7584
rect 38666 7648 38982 7649
rect 38666 7584 38672 7648
rect 38736 7584 38752 7648
rect 38816 7584 38832 7648
rect 38896 7584 38912 7648
rect 38976 7584 38982 7648
rect 38666 7583 38982 7584
rect 5661 7104 5977 7105
rect 5661 7040 5667 7104
rect 5731 7040 5747 7104
rect 5811 7040 5827 7104
rect 5891 7040 5907 7104
rect 5971 7040 5977 7104
rect 5661 7039 5977 7040
rect 15091 7104 15407 7105
rect 15091 7040 15097 7104
rect 15161 7040 15177 7104
rect 15241 7040 15257 7104
rect 15321 7040 15337 7104
rect 15401 7040 15407 7104
rect 15091 7039 15407 7040
rect 24521 7104 24837 7105
rect 24521 7040 24527 7104
rect 24591 7040 24607 7104
rect 24671 7040 24687 7104
rect 24751 7040 24767 7104
rect 24831 7040 24837 7104
rect 24521 7039 24837 7040
rect 33951 7104 34267 7105
rect 33951 7040 33957 7104
rect 34021 7040 34037 7104
rect 34101 7040 34117 7104
rect 34181 7040 34197 7104
rect 34261 7040 34267 7104
rect 33951 7039 34267 7040
rect 10376 6560 10692 6561
rect 10376 6496 10382 6560
rect 10446 6496 10462 6560
rect 10526 6496 10542 6560
rect 10606 6496 10622 6560
rect 10686 6496 10692 6560
rect 10376 6495 10692 6496
rect 19806 6560 20122 6561
rect 19806 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20052 6560
rect 20116 6496 20122 6560
rect 19806 6495 20122 6496
rect 29236 6560 29552 6561
rect 29236 6496 29242 6560
rect 29306 6496 29322 6560
rect 29386 6496 29402 6560
rect 29466 6496 29482 6560
rect 29546 6496 29552 6560
rect 29236 6495 29552 6496
rect 38666 6560 38982 6561
rect 38666 6496 38672 6560
rect 38736 6496 38752 6560
rect 38816 6496 38832 6560
rect 38896 6496 38912 6560
rect 38976 6496 38982 6560
rect 38666 6495 38982 6496
rect 38469 6218 38535 6221
rect 39200 6218 40000 6248
rect 38469 6216 40000 6218
rect 38469 6160 38474 6216
rect 38530 6160 40000 6216
rect 38469 6158 40000 6160
rect 38469 6155 38535 6158
rect 39200 6128 40000 6158
rect 5661 6016 5977 6017
rect 5661 5952 5667 6016
rect 5731 5952 5747 6016
rect 5811 5952 5827 6016
rect 5891 5952 5907 6016
rect 5971 5952 5977 6016
rect 5661 5951 5977 5952
rect 15091 6016 15407 6017
rect 15091 5952 15097 6016
rect 15161 5952 15177 6016
rect 15241 5952 15257 6016
rect 15321 5952 15337 6016
rect 15401 5952 15407 6016
rect 15091 5951 15407 5952
rect 24521 6016 24837 6017
rect 24521 5952 24527 6016
rect 24591 5952 24607 6016
rect 24671 5952 24687 6016
rect 24751 5952 24767 6016
rect 24831 5952 24837 6016
rect 24521 5951 24837 5952
rect 33951 6016 34267 6017
rect 33951 5952 33957 6016
rect 34021 5952 34037 6016
rect 34101 5952 34117 6016
rect 34181 5952 34197 6016
rect 34261 5952 34267 6016
rect 33951 5951 34267 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 10376 5472 10692 5473
rect 10376 5408 10382 5472
rect 10446 5408 10462 5472
rect 10526 5408 10542 5472
rect 10606 5408 10622 5472
rect 10686 5408 10692 5472
rect 10376 5407 10692 5408
rect 19806 5472 20122 5473
rect 19806 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20052 5472
rect 20116 5408 20122 5472
rect 19806 5407 20122 5408
rect 29236 5472 29552 5473
rect 29236 5408 29242 5472
rect 29306 5408 29322 5472
rect 29386 5408 29402 5472
rect 29466 5408 29482 5472
rect 29546 5408 29552 5472
rect 29236 5407 29552 5408
rect 38666 5472 38982 5473
rect 38666 5408 38672 5472
rect 38736 5408 38752 5472
rect 38816 5408 38832 5472
rect 38896 5408 38912 5472
rect 38976 5408 38982 5472
rect 38666 5407 38982 5408
rect 5661 4928 5977 4929
rect 5661 4864 5667 4928
rect 5731 4864 5747 4928
rect 5811 4864 5827 4928
rect 5891 4864 5907 4928
rect 5971 4864 5977 4928
rect 5661 4863 5977 4864
rect 15091 4928 15407 4929
rect 15091 4864 15097 4928
rect 15161 4864 15177 4928
rect 15241 4864 15257 4928
rect 15321 4864 15337 4928
rect 15401 4864 15407 4928
rect 15091 4863 15407 4864
rect 24521 4928 24837 4929
rect 24521 4864 24527 4928
rect 24591 4864 24607 4928
rect 24671 4864 24687 4928
rect 24751 4864 24767 4928
rect 24831 4864 24837 4928
rect 24521 4863 24837 4864
rect 33951 4928 34267 4929
rect 33951 4864 33957 4928
rect 34021 4864 34037 4928
rect 34101 4864 34117 4928
rect 34181 4864 34197 4928
rect 34261 4864 34267 4928
rect 33951 4863 34267 4864
rect 10376 4384 10692 4385
rect 10376 4320 10382 4384
rect 10446 4320 10462 4384
rect 10526 4320 10542 4384
rect 10606 4320 10622 4384
rect 10686 4320 10692 4384
rect 10376 4319 10692 4320
rect 19806 4384 20122 4385
rect 19806 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20052 4384
rect 20116 4320 20122 4384
rect 19806 4319 20122 4320
rect 29236 4384 29552 4385
rect 29236 4320 29242 4384
rect 29306 4320 29322 4384
rect 29386 4320 29402 4384
rect 29466 4320 29482 4384
rect 29546 4320 29552 4384
rect 29236 4319 29552 4320
rect 38666 4384 38982 4385
rect 38666 4320 38672 4384
rect 38736 4320 38752 4384
rect 38816 4320 38832 4384
rect 38896 4320 38912 4384
rect 38976 4320 38982 4384
rect 38666 4319 38982 4320
rect 5661 3840 5977 3841
rect 5661 3776 5667 3840
rect 5731 3776 5747 3840
rect 5811 3776 5827 3840
rect 5891 3776 5907 3840
rect 5971 3776 5977 3840
rect 5661 3775 5977 3776
rect 15091 3840 15407 3841
rect 15091 3776 15097 3840
rect 15161 3776 15177 3840
rect 15241 3776 15257 3840
rect 15321 3776 15337 3840
rect 15401 3776 15407 3840
rect 15091 3775 15407 3776
rect 24521 3840 24837 3841
rect 24521 3776 24527 3840
rect 24591 3776 24607 3840
rect 24671 3776 24687 3840
rect 24751 3776 24767 3840
rect 24831 3776 24837 3840
rect 24521 3775 24837 3776
rect 33951 3840 34267 3841
rect 33951 3776 33957 3840
rect 34021 3776 34037 3840
rect 34101 3776 34117 3840
rect 34181 3776 34197 3840
rect 34261 3776 34267 3840
rect 33951 3775 34267 3776
rect 38469 3498 38535 3501
rect 39200 3498 40000 3528
rect 38469 3496 40000 3498
rect 38469 3440 38474 3496
rect 38530 3440 40000 3496
rect 38469 3438 40000 3440
rect 38469 3435 38535 3438
rect 39200 3408 40000 3438
rect 10376 3296 10692 3297
rect 10376 3232 10382 3296
rect 10446 3232 10462 3296
rect 10526 3232 10542 3296
rect 10606 3232 10622 3296
rect 10686 3232 10692 3296
rect 10376 3231 10692 3232
rect 19806 3296 20122 3297
rect 19806 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20052 3296
rect 20116 3232 20122 3296
rect 19806 3231 20122 3232
rect 29236 3296 29552 3297
rect 29236 3232 29242 3296
rect 29306 3232 29322 3296
rect 29386 3232 29402 3296
rect 29466 3232 29482 3296
rect 29546 3232 29552 3296
rect 29236 3231 29552 3232
rect 38666 3296 38982 3297
rect 38666 3232 38672 3296
rect 38736 3232 38752 3296
rect 38816 3232 38832 3296
rect 38896 3232 38912 3296
rect 38976 3232 38982 3296
rect 38666 3231 38982 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 5661 2752 5977 2753
rect 5661 2688 5667 2752
rect 5731 2688 5747 2752
rect 5811 2688 5827 2752
rect 5891 2688 5907 2752
rect 5971 2688 5977 2752
rect 5661 2687 5977 2688
rect 15091 2752 15407 2753
rect 15091 2688 15097 2752
rect 15161 2688 15177 2752
rect 15241 2688 15257 2752
rect 15321 2688 15337 2752
rect 15401 2688 15407 2752
rect 15091 2687 15407 2688
rect 24521 2752 24837 2753
rect 24521 2688 24527 2752
rect 24591 2688 24607 2752
rect 24671 2688 24687 2752
rect 24751 2688 24767 2752
rect 24831 2688 24837 2752
rect 24521 2687 24837 2688
rect 33951 2752 34267 2753
rect 33951 2688 33957 2752
rect 34021 2688 34037 2752
rect 34101 2688 34117 2752
rect 34181 2688 34197 2752
rect 34261 2688 34267 2752
rect 33951 2687 34267 2688
rect 10376 2208 10692 2209
rect 10376 2144 10382 2208
rect 10446 2144 10462 2208
rect 10526 2144 10542 2208
rect 10606 2144 10622 2208
rect 10686 2144 10692 2208
rect 10376 2143 10692 2144
rect 19806 2208 20122 2209
rect 19806 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20052 2208
rect 20116 2144 20122 2208
rect 19806 2143 20122 2144
rect 29236 2208 29552 2209
rect 29236 2144 29242 2208
rect 29306 2144 29322 2208
rect 29386 2144 29402 2208
rect 29466 2144 29482 2208
rect 29546 2144 29552 2208
rect 29236 2143 29552 2144
rect 38666 2208 38982 2209
rect 38666 2144 38672 2208
rect 38736 2144 38752 2208
rect 38816 2144 38832 2208
rect 38896 2144 38912 2208
rect 38976 2144 38982 2208
rect 38666 2143 38982 2144
rect 38469 778 38535 781
rect 39200 778 40000 808
rect 38469 776 40000 778
rect 38469 720 38474 776
rect 38530 720 40000 776
rect 38469 718 40000 720
rect 38469 715 38535 718
rect 39200 688 40000 718
<< via3 >>
rect 10382 9820 10446 9824
rect 10382 9764 10386 9820
rect 10386 9764 10442 9820
rect 10442 9764 10446 9820
rect 10382 9760 10446 9764
rect 10462 9820 10526 9824
rect 10462 9764 10466 9820
rect 10466 9764 10522 9820
rect 10522 9764 10526 9820
rect 10462 9760 10526 9764
rect 10542 9820 10606 9824
rect 10542 9764 10546 9820
rect 10546 9764 10602 9820
rect 10602 9764 10606 9820
rect 10542 9760 10606 9764
rect 10622 9820 10686 9824
rect 10622 9764 10626 9820
rect 10626 9764 10682 9820
rect 10682 9764 10686 9820
rect 10622 9760 10686 9764
rect 19812 9820 19876 9824
rect 19812 9764 19816 9820
rect 19816 9764 19872 9820
rect 19872 9764 19876 9820
rect 19812 9760 19876 9764
rect 19892 9820 19956 9824
rect 19892 9764 19896 9820
rect 19896 9764 19952 9820
rect 19952 9764 19956 9820
rect 19892 9760 19956 9764
rect 19972 9820 20036 9824
rect 19972 9764 19976 9820
rect 19976 9764 20032 9820
rect 20032 9764 20036 9820
rect 19972 9760 20036 9764
rect 20052 9820 20116 9824
rect 20052 9764 20056 9820
rect 20056 9764 20112 9820
rect 20112 9764 20116 9820
rect 20052 9760 20116 9764
rect 29242 9820 29306 9824
rect 29242 9764 29246 9820
rect 29246 9764 29302 9820
rect 29302 9764 29306 9820
rect 29242 9760 29306 9764
rect 29322 9820 29386 9824
rect 29322 9764 29326 9820
rect 29326 9764 29382 9820
rect 29382 9764 29386 9820
rect 29322 9760 29386 9764
rect 29402 9820 29466 9824
rect 29402 9764 29406 9820
rect 29406 9764 29462 9820
rect 29462 9764 29466 9820
rect 29402 9760 29466 9764
rect 29482 9820 29546 9824
rect 29482 9764 29486 9820
rect 29486 9764 29542 9820
rect 29542 9764 29546 9820
rect 29482 9760 29546 9764
rect 38672 9820 38736 9824
rect 38672 9764 38676 9820
rect 38676 9764 38732 9820
rect 38732 9764 38736 9820
rect 38672 9760 38736 9764
rect 38752 9820 38816 9824
rect 38752 9764 38756 9820
rect 38756 9764 38812 9820
rect 38812 9764 38816 9820
rect 38752 9760 38816 9764
rect 38832 9820 38896 9824
rect 38832 9764 38836 9820
rect 38836 9764 38892 9820
rect 38892 9764 38896 9820
rect 38832 9760 38896 9764
rect 38912 9820 38976 9824
rect 38912 9764 38916 9820
rect 38916 9764 38972 9820
rect 38972 9764 38976 9820
rect 38912 9760 38976 9764
rect 5667 9276 5731 9280
rect 5667 9220 5671 9276
rect 5671 9220 5727 9276
rect 5727 9220 5731 9276
rect 5667 9216 5731 9220
rect 5747 9276 5811 9280
rect 5747 9220 5751 9276
rect 5751 9220 5807 9276
rect 5807 9220 5811 9276
rect 5747 9216 5811 9220
rect 5827 9276 5891 9280
rect 5827 9220 5831 9276
rect 5831 9220 5887 9276
rect 5887 9220 5891 9276
rect 5827 9216 5891 9220
rect 5907 9276 5971 9280
rect 5907 9220 5911 9276
rect 5911 9220 5967 9276
rect 5967 9220 5971 9276
rect 5907 9216 5971 9220
rect 15097 9276 15161 9280
rect 15097 9220 15101 9276
rect 15101 9220 15157 9276
rect 15157 9220 15161 9276
rect 15097 9216 15161 9220
rect 15177 9276 15241 9280
rect 15177 9220 15181 9276
rect 15181 9220 15237 9276
rect 15237 9220 15241 9276
rect 15177 9216 15241 9220
rect 15257 9276 15321 9280
rect 15257 9220 15261 9276
rect 15261 9220 15317 9276
rect 15317 9220 15321 9276
rect 15257 9216 15321 9220
rect 15337 9276 15401 9280
rect 15337 9220 15341 9276
rect 15341 9220 15397 9276
rect 15397 9220 15401 9276
rect 15337 9216 15401 9220
rect 24527 9276 24591 9280
rect 24527 9220 24531 9276
rect 24531 9220 24587 9276
rect 24587 9220 24591 9276
rect 24527 9216 24591 9220
rect 24607 9276 24671 9280
rect 24607 9220 24611 9276
rect 24611 9220 24667 9276
rect 24667 9220 24671 9276
rect 24607 9216 24671 9220
rect 24687 9276 24751 9280
rect 24687 9220 24691 9276
rect 24691 9220 24747 9276
rect 24747 9220 24751 9276
rect 24687 9216 24751 9220
rect 24767 9276 24831 9280
rect 24767 9220 24771 9276
rect 24771 9220 24827 9276
rect 24827 9220 24831 9276
rect 24767 9216 24831 9220
rect 33957 9276 34021 9280
rect 33957 9220 33961 9276
rect 33961 9220 34017 9276
rect 34017 9220 34021 9276
rect 33957 9216 34021 9220
rect 34037 9276 34101 9280
rect 34037 9220 34041 9276
rect 34041 9220 34097 9276
rect 34097 9220 34101 9276
rect 34037 9216 34101 9220
rect 34117 9276 34181 9280
rect 34117 9220 34121 9276
rect 34121 9220 34177 9276
rect 34177 9220 34181 9276
rect 34117 9216 34181 9220
rect 34197 9276 34261 9280
rect 34197 9220 34201 9276
rect 34201 9220 34257 9276
rect 34257 9220 34261 9276
rect 34197 9216 34261 9220
rect 10382 8732 10446 8736
rect 10382 8676 10386 8732
rect 10386 8676 10442 8732
rect 10442 8676 10446 8732
rect 10382 8672 10446 8676
rect 10462 8732 10526 8736
rect 10462 8676 10466 8732
rect 10466 8676 10522 8732
rect 10522 8676 10526 8732
rect 10462 8672 10526 8676
rect 10542 8732 10606 8736
rect 10542 8676 10546 8732
rect 10546 8676 10602 8732
rect 10602 8676 10606 8732
rect 10542 8672 10606 8676
rect 10622 8732 10686 8736
rect 10622 8676 10626 8732
rect 10626 8676 10682 8732
rect 10682 8676 10686 8732
rect 10622 8672 10686 8676
rect 19812 8732 19876 8736
rect 19812 8676 19816 8732
rect 19816 8676 19872 8732
rect 19872 8676 19876 8732
rect 19812 8672 19876 8676
rect 19892 8732 19956 8736
rect 19892 8676 19896 8732
rect 19896 8676 19952 8732
rect 19952 8676 19956 8732
rect 19892 8672 19956 8676
rect 19972 8732 20036 8736
rect 19972 8676 19976 8732
rect 19976 8676 20032 8732
rect 20032 8676 20036 8732
rect 19972 8672 20036 8676
rect 20052 8732 20116 8736
rect 20052 8676 20056 8732
rect 20056 8676 20112 8732
rect 20112 8676 20116 8732
rect 20052 8672 20116 8676
rect 29242 8732 29306 8736
rect 29242 8676 29246 8732
rect 29246 8676 29302 8732
rect 29302 8676 29306 8732
rect 29242 8672 29306 8676
rect 29322 8732 29386 8736
rect 29322 8676 29326 8732
rect 29326 8676 29382 8732
rect 29382 8676 29386 8732
rect 29322 8672 29386 8676
rect 29402 8732 29466 8736
rect 29402 8676 29406 8732
rect 29406 8676 29462 8732
rect 29462 8676 29466 8732
rect 29402 8672 29466 8676
rect 29482 8732 29546 8736
rect 29482 8676 29486 8732
rect 29486 8676 29542 8732
rect 29542 8676 29546 8732
rect 29482 8672 29546 8676
rect 38672 8732 38736 8736
rect 38672 8676 38676 8732
rect 38676 8676 38732 8732
rect 38732 8676 38736 8732
rect 38672 8672 38736 8676
rect 38752 8732 38816 8736
rect 38752 8676 38756 8732
rect 38756 8676 38812 8732
rect 38812 8676 38816 8732
rect 38752 8672 38816 8676
rect 38832 8732 38896 8736
rect 38832 8676 38836 8732
rect 38836 8676 38892 8732
rect 38892 8676 38896 8732
rect 38832 8672 38896 8676
rect 38912 8732 38976 8736
rect 38912 8676 38916 8732
rect 38916 8676 38972 8732
rect 38972 8676 38976 8732
rect 38912 8672 38976 8676
rect 5667 8188 5731 8192
rect 5667 8132 5671 8188
rect 5671 8132 5727 8188
rect 5727 8132 5731 8188
rect 5667 8128 5731 8132
rect 5747 8188 5811 8192
rect 5747 8132 5751 8188
rect 5751 8132 5807 8188
rect 5807 8132 5811 8188
rect 5747 8128 5811 8132
rect 5827 8188 5891 8192
rect 5827 8132 5831 8188
rect 5831 8132 5887 8188
rect 5887 8132 5891 8188
rect 5827 8128 5891 8132
rect 5907 8188 5971 8192
rect 5907 8132 5911 8188
rect 5911 8132 5967 8188
rect 5967 8132 5971 8188
rect 5907 8128 5971 8132
rect 15097 8188 15161 8192
rect 15097 8132 15101 8188
rect 15101 8132 15157 8188
rect 15157 8132 15161 8188
rect 15097 8128 15161 8132
rect 15177 8188 15241 8192
rect 15177 8132 15181 8188
rect 15181 8132 15237 8188
rect 15237 8132 15241 8188
rect 15177 8128 15241 8132
rect 15257 8188 15321 8192
rect 15257 8132 15261 8188
rect 15261 8132 15317 8188
rect 15317 8132 15321 8188
rect 15257 8128 15321 8132
rect 15337 8188 15401 8192
rect 15337 8132 15341 8188
rect 15341 8132 15397 8188
rect 15397 8132 15401 8188
rect 15337 8128 15401 8132
rect 24527 8188 24591 8192
rect 24527 8132 24531 8188
rect 24531 8132 24587 8188
rect 24587 8132 24591 8188
rect 24527 8128 24591 8132
rect 24607 8188 24671 8192
rect 24607 8132 24611 8188
rect 24611 8132 24667 8188
rect 24667 8132 24671 8188
rect 24607 8128 24671 8132
rect 24687 8188 24751 8192
rect 24687 8132 24691 8188
rect 24691 8132 24747 8188
rect 24747 8132 24751 8188
rect 24687 8128 24751 8132
rect 24767 8188 24831 8192
rect 24767 8132 24771 8188
rect 24771 8132 24827 8188
rect 24827 8132 24831 8188
rect 24767 8128 24831 8132
rect 33957 8188 34021 8192
rect 33957 8132 33961 8188
rect 33961 8132 34017 8188
rect 34017 8132 34021 8188
rect 33957 8128 34021 8132
rect 34037 8188 34101 8192
rect 34037 8132 34041 8188
rect 34041 8132 34097 8188
rect 34097 8132 34101 8188
rect 34037 8128 34101 8132
rect 34117 8188 34181 8192
rect 34117 8132 34121 8188
rect 34121 8132 34177 8188
rect 34177 8132 34181 8188
rect 34117 8128 34181 8132
rect 34197 8188 34261 8192
rect 34197 8132 34201 8188
rect 34201 8132 34257 8188
rect 34257 8132 34261 8188
rect 34197 8128 34261 8132
rect 10382 7644 10446 7648
rect 10382 7588 10386 7644
rect 10386 7588 10442 7644
rect 10442 7588 10446 7644
rect 10382 7584 10446 7588
rect 10462 7644 10526 7648
rect 10462 7588 10466 7644
rect 10466 7588 10522 7644
rect 10522 7588 10526 7644
rect 10462 7584 10526 7588
rect 10542 7644 10606 7648
rect 10542 7588 10546 7644
rect 10546 7588 10602 7644
rect 10602 7588 10606 7644
rect 10542 7584 10606 7588
rect 10622 7644 10686 7648
rect 10622 7588 10626 7644
rect 10626 7588 10682 7644
rect 10682 7588 10686 7644
rect 10622 7584 10686 7588
rect 19812 7644 19876 7648
rect 19812 7588 19816 7644
rect 19816 7588 19872 7644
rect 19872 7588 19876 7644
rect 19812 7584 19876 7588
rect 19892 7644 19956 7648
rect 19892 7588 19896 7644
rect 19896 7588 19952 7644
rect 19952 7588 19956 7644
rect 19892 7584 19956 7588
rect 19972 7644 20036 7648
rect 19972 7588 19976 7644
rect 19976 7588 20032 7644
rect 20032 7588 20036 7644
rect 19972 7584 20036 7588
rect 20052 7644 20116 7648
rect 20052 7588 20056 7644
rect 20056 7588 20112 7644
rect 20112 7588 20116 7644
rect 20052 7584 20116 7588
rect 29242 7644 29306 7648
rect 29242 7588 29246 7644
rect 29246 7588 29302 7644
rect 29302 7588 29306 7644
rect 29242 7584 29306 7588
rect 29322 7644 29386 7648
rect 29322 7588 29326 7644
rect 29326 7588 29382 7644
rect 29382 7588 29386 7644
rect 29322 7584 29386 7588
rect 29402 7644 29466 7648
rect 29402 7588 29406 7644
rect 29406 7588 29462 7644
rect 29462 7588 29466 7644
rect 29402 7584 29466 7588
rect 29482 7644 29546 7648
rect 29482 7588 29486 7644
rect 29486 7588 29542 7644
rect 29542 7588 29546 7644
rect 29482 7584 29546 7588
rect 38672 7644 38736 7648
rect 38672 7588 38676 7644
rect 38676 7588 38732 7644
rect 38732 7588 38736 7644
rect 38672 7584 38736 7588
rect 38752 7644 38816 7648
rect 38752 7588 38756 7644
rect 38756 7588 38812 7644
rect 38812 7588 38816 7644
rect 38752 7584 38816 7588
rect 38832 7644 38896 7648
rect 38832 7588 38836 7644
rect 38836 7588 38892 7644
rect 38892 7588 38896 7644
rect 38832 7584 38896 7588
rect 38912 7644 38976 7648
rect 38912 7588 38916 7644
rect 38916 7588 38972 7644
rect 38972 7588 38976 7644
rect 38912 7584 38976 7588
rect 5667 7100 5731 7104
rect 5667 7044 5671 7100
rect 5671 7044 5727 7100
rect 5727 7044 5731 7100
rect 5667 7040 5731 7044
rect 5747 7100 5811 7104
rect 5747 7044 5751 7100
rect 5751 7044 5807 7100
rect 5807 7044 5811 7100
rect 5747 7040 5811 7044
rect 5827 7100 5891 7104
rect 5827 7044 5831 7100
rect 5831 7044 5887 7100
rect 5887 7044 5891 7100
rect 5827 7040 5891 7044
rect 5907 7100 5971 7104
rect 5907 7044 5911 7100
rect 5911 7044 5967 7100
rect 5967 7044 5971 7100
rect 5907 7040 5971 7044
rect 15097 7100 15161 7104
rect 15097 7044 15101 7100
rect 15101 7044 15157 7100
rect 15157 7044 15161 7100
rect 15097 7040 15161 7044
rect 15177 7100 15241 7104
rect 15177 7044 15181 7100
rect 15181 7044 15237 7100
rect 15237 7044 15241 7100
rect 15177 7040 15241 7044
rect 15257 7100 15321 7104
rect 15257 7044 15261 7100
rect 15261 7044 15317 7100
rect 15317 7044 15321 7100
rect 15257 7040 15321 7044
rect 15337 7100 15401 7104
rect 15337 7044 15341 7100
rect 15341 7044 15397 7100
rect 15397 7044 15401 7100
rect 15337 7040 15401 7044
rect 24527 7100 24591 7104
rect 24527 7044 24531 7100
rect 24531 7044 24587 7100
rect 24587 7044 24591 7100
rect 24527 7040 24591 7044
rect 24607 7100 24671 7104
rect 24607 7044 24611 7100
rect 24611 7044 24667 7100
rect 24667 7044 24671 7100
rect 24607 7040 24671 7044
rect 24687 7100 24751 7104
rect 24687 7044 24691 7100
rect 24691 7044 24747 7100
rect 24747 7044 24751 7100
rect 24687 7040 24751 7044
rect 24767 7100 24831 7104
rect 24767 7044 24771 7100
rect 24771 7044 24827 7100
rect 24827 7044 24831 7100
rect 24767 7040 24831 7044
rect 33957 7100 34021 7104
rect 33957 7044 33961 7100
rect 33961 7044 34017 7100
rect 34017 7044 34021 7100
rect 33957 7040 34021 7044
rect 34037 7100 34101 7104
rect 34037 7044 34041 7100
rect 34041 7044 34097 7100
rect 34097 7044 34101 7100
rect 34037 7040 34101 7044
rect 34117 7100 34181 7104
rect 34117 7044 34121 7100
rect 34121 7044 34177 7100
rect 34177 7044 34181 7100
rect 34117 7040 34181 7044
rect 34197 7100 34261 7104
rect 34197 7044 34201 7100
rect 34201 7044 34257 7100
rect 34257 7044 34261 7100
rect 34197 7040 34261 7044
rect 10382 6556 10446 6560
rect 10382 6500 10386 6556
rect 10386 6500 10442 6556
rect 10442 6500 10446 6556
rect 10382 6496 10446 6500
rect 10462 6556 10526 6560
rect 10462 6500 10466 6556
rect 10466 6500 10522 6556
rect 10522 6500 10526 6556
rect 10462 6496 10526 6500
rect 10542 6556 10606 6560
rect 10542 6500 10546 6556
rect 10546 6500 10602 6556
rect 10602 6500 10606 6556
rect 10542 6496 10606 6500
rect 10622 6556 10686 6560
rect 10622 6500 10626 6556
rect 10626 6500 10682 6556
rect 10682 6500 10686 6556
rect 10622 6496 10686 6500
rect 19812 6556 19876 6560
rect 19812 6500 19816 6556
rect 19816 6500 19872 6556
rect 19872 6500 19876 6556
rect 19812 6496 19876 6500
rect 19892 6556 19956 6560
rect 19892 6500 19896 6556
rect 19896 6500 19952 6556
rect 19952 6500 19956 6556
rect 19892 6496 19956 6500
rect 19972 6556 20036 6560
rect 19972 6500 19976 6556
rect 19976 6500 20032 6556
rect 20032 6500 20036 6556
rect 19972 6496 20036 6500
rect 20052 6556 20116 6560
rect 20052 6500 20056 6556
rect 20056 6500 20112 6556
rect 20112 6500 20116 6556
rect 20052 6496 20116 6500
rect 29242 6556 29306 6560
rect 29242 6500 29246 6556
rect 29246 6500 29302 6556
rect 29302 6500 29306 6556
rect 29242 6496 29306 6500
rect 29322 6556 29386 6560
rect 29322 6500 29326 6556
rect 29326 6500 29382 6556
rect 29382 6500 29386 6556
rect 29322 6496 29386 6500
rect 29402 6556 29466 6560
rect 29402 6500 29406 6556
rect 29406 6500 29462 6556
rect 29462 6500 29466 6556
rect 29402 6496 29466 6500
rect 29482 6556 29546 6560
rect 29482 6500 29486 6556
rect 29486 6500 29542 6556
rect 29542 6500 29546 6556
rect 29482 6496 29546 6500
rect 38672 6556 38736 6560
rect 38672 6500 38676 6556
rect 38676 6500 38732 6556
rect 38732 6500 38736 6556
rect 38672 6496 38736 6500
rect 38752 6556 38816 6560
rect 38752 6500 38756 6556
rect 38756 6500 38812 6556
rect 38812 6500 38816 6556
rect 38752 6496 38816 6500
rect 38832 6556 38896 6560
rect 38832 6500 38836 6556
rect 38836 6500 38892 6556
rect 38892 6500 38896 6556
rect 38832 6496 38896 6500
rect 38912 6556 38976 6560
rect 38912 6500 38916 6556
rect 38916 6500 38972 6556
rect 38972 6500 38976 6556
rect 38912 6496 38976 6500
rect 5667 6012 5731 6016
rect 5667 5956 5671 6012
rect 5671 5956 5727 6012
rect 5727 5956 5731 6012
rect 5667 5952 5731 5956
rect 5747 6012 5811 6016
rect 5747 5956 5751 6012
rect 5751 5956 5807 6012
rect 5807 5956 5811 6012
rect 5747 5952 5811 5956
rect 5827 6012 5891 6016
rect 5827 5956 5831 6012
rect 5831 5956 5887 6012
rect 5887 5956 5891 6012
rect 5827 5952 5891 5956
rect 5907 6012 5971 6016
rect 5907 5956 5911 6012
rect 5911 5956 5967 6012
rect 5967 5956 5971 6012
rect 5907 5952 5971 5956
rect 15097 6012 15161 6016
rect 15097 5956 15101 6012
rect 15101 5956 15157 6012
rect 15157 5956 15161 6012
rect 15097 5952 15161 5956
rect 15177 6012 15241 6016
rect 15177 5956 15181 6012
rect 15181 5956 15237 6012
rect 15237 5956 15241 6012
rect 15177 5952 15241 5956
rect 15257 6012 15321 6016
rect 15257 5956 15261 6012
rect 15261 5956 15317 6012
rect 15317 5956 15321 6012
rect 15257 5952 15321 5956
rect 15337 6012 15401 6016
rect 15337 5956 15341 6012
rect 15341 5956 15397 6012
rect 15397 5956 15401 6012
rect 15337 5952 15401 5956
rect 24527 6012 24591 6016
rect 24527 5956 24531 6012
rect 24531 5956 24587 6012
rect 24587 5956 24591 6012
rect 24527 5952 24591 5956
rect 24607 6012 24671 6016
rect 24607 5956 24611 6012
rect 24611 5956 24667 6012
rect 24667 5956 24671 6012
rect 24607 5952 24671 5956
rect 24687 6012 24751 6016
rect 24687 5956 24691 6012
rect 24691 5956 24747 6012
rect 24747 5956 24751 6012
rect 24687 5952 24751 5956
rect 24767 6012 24831 6016
rect 24767 5956 24771 6012
rect 24771 5956 24827 6012
rect 24827 5956 24831 6012
rect 24767 5952 24831 5956
rect 33957 6012 34021 6016
rect 33957 5956 33961 6012
rect 33961 5956 34017 6012
rect 34017 5956 34021 6012
rect 33957 5952 34021 5956
rect 34037 6012 34101 6016
rect 34037 5956 34041 6012
rect 34041 5956 34097 6012
rect 34097 5956 34101 6012
rect 34037 5952 34101 5956
rect 34117 6012 34181 6016
rect 34117 5956 34121 6012
rect 34121 5956 34177 6012
rect 34177 5956 34181 6012
rect 34117 5952 34181 5956
rect 34197 6012 34261 6016
rect 34197 5956 34201 6012
rect 34201 5956 34257 6012
rect 34257 5956 34261 6012
rect 34197 5952 34261 5956
rect 10382 5468 10446 5472
rect 10382 5412 10386 5468
rect 10386 5412 10442 5468
rect 10442 5412 10446 5468
rect 10382 5408 10446 5412
rect 10462 5468 10526 5472
rect 10462 5412 10466 5468
rect 10466 5412 10522 5468
rect 10522 5412 10526 5468
rect 10462 5408 10526 5412
rect 10542 5468 10606 5472
rect 10542 5412 10546 5468
rect 10546 5412 10602 5468
rect 10602 5412 10606 5468
rect 10542 5408 10606 5412
rect 10622 5468 10686 5472
rect 10622 5412 10626 5468
rect 10626 5412 10682 5468
rect 10682 5412 10686 5468
rect 10622 5408 10686 5412
rect 19812 5468 19876 5472
rect 19812 5412 19816 5468
rect 19816 5412 19872 5468
rect 19872 5412 19876 5468
rect 19812 5408 19876 5412
rect 19892 5468 19956 5472
rect 19892 5412 19896 5468
rect 19896 5412 19952 5468
rect 19952 5412 19956 5468
rect 19892 5408 19956 5412
rect 19972 5468 20036 5472
rect 19972 5412 19976 5468
rect 19976 5412 20032 5468
rect 20032 5412 20036 5468
rect 19972 5408 20036 5412
rect 20052 5468 20116 5472
rect 20052 5412 20056 5468
rect 20056 5412 20112 5468
rect 20112 5412 20116 5468
rect 20052 5408 20116 5412
rect 29242 5468 29306 5472
rect 29242 5412 29246 5468
rect 29246 5412 29302 5468
rect 29302 5412 29306 5468
rect 29242 5408 29306 5412
rect 29322 5468 29386 5472
rect 29322 5412 29326 5468
rect 29326 5412 29382 5468
rect 29382 5412 29386 5468
rect 29322 5408 29386 5412
rect 29402 5468 29466 5472
rect 29402 5412 29406 5468
rect 29406 5412 29462 5468
rect 29462 5412 29466 5468
rect 29402 5408 29466 5412
rect 29482 5468 29546 5472
rect 29482 5412 29486 5468
rect 29486 5412 29542 5468
rect 29542 5412 29546 5468
rect 29482 5408 29546 5412
rect 38672 5468 38736 5472
rect 38672 5412 38676 5468
rect 38676 5412 38732 5468
rect 38732 5412 38736 5468
rect 38672 5408 38736 5412
rect 38752 5468 38816 5472
rect 38752 5412 38756 5468
rect 38756 5412 38812 5468
rect 38812 5412 38816 5468
rect 38752 5408 38816 5412
rect 38832 5468 38896 5472
rect 38832 5412 38836 5468
rect 38836 5412 38892 5468
rect 38892 5412 38896 5468
rect 38832 5408 38896 5412
rect 38912 5468 38976 5472
rect 38912 5412 38916 5468
rect 38916 5412 38972 5468
rect 38972 5412 38976 5468
rect 38912 5408 38976 5412
rect 5667 4924 5731 4928
rect 5667 4868 5671 4924
rect 5671 4868 5727 4924
rect 5727 4868 5731 4924
rect 5667 4864 5731 4868
rect 5747 4924 5811 4928
rect 5747 4868 5751 4924
rect 5751 4868 5807 4924
rect 5807 4868 5811 4924
rect 5747 4864 5811 4868
rect 5827 4924 5891 4928
rect 5827 4868 5831 4924
rect 5831 4868 5887 4924
rect 5887 4868 5891 4924
rect 5827 4864 5891 4868
rect 5907 4924 5971 4928
rect 5907 4868 5911 4924
rect 5911 4868 5967 4924
rect 5967 4868 5971 4924
rect 5907 4864 5971 4868
rect 15097 4924 15161 4928
rect 15097 4868 15101 4924
rect 15101 4868 15157 4924
rect 15157 4868 15161 4924
rect 15097 4864 15161 4868
rect 15177 4924 15241 4928
rect 15177 4868 15181 4924
rect 15181 4868 15237 4924
rect 15237 4868 15241 4924
rect 15177 4864 15241 4868
rect 15257 4924 15321 4928
rect 15257 4868 15261 4924
rect 15261 4868 15317 4924
rect 15317 4868 15321 4924
rect 15257 4864 15321 4868
rect 15337 4924 15401 4928
rect 15337 4868 15341 4924
rect 15341 4868 15397 4924
rect 15397 4868 15401 4924
rect 15337 4864 15401 4868
rect 24527 4924 24591 4928
rect 24527 4868 24531 4924
rect 24531 4868 24587 4924
rect 24587 4868 24591 4924
rect 24527 4864 24591 4868
rect 24607 4924 24671 4928
rect 24607 4868 24611 4924
rect 24611 4868 24667 4924
rect 24667 4868 24671 4924
rect 24607 4864 24671 4868
rect 24687 4924 24751 4928
rect 24687 4868 24691 4924
rect 24691 4868 24747 4924
rect 24747 4868 24751 4924
rect 24687 4864 24751 4868
rect 24767 4924 24831 4928
rect 24767 4868 24771 4924
rect 24771 4868 24827 4924
rect 24827 4868 24831 4924
rect 24767 4864 24831 4868
rect 33957 4924 34021 4928
rect 33957 4868 33961 4924
rect 33961 4868 34017 4924
rect 34017 4868 34021 4924
rect 33957 4864 34021 4868
rect 34037 4924 34101 4928
rect 34037 4868 34041 4924
rect 34041 4868 34097 4924
rect 34097 4868 34101 4924
rect 34037 4864 34101 4868
rect 34117 4924 34181 4928
rect 34117 4868 34121 4924
rect 34121 4868 34177 4924
rect 34177 4868 34181 4924
rect 34117 4864 34181 4868
rect 34197 4924 34261 4928
rect 34197 4868 34201 4924
rect 34201 4868 34257 4924
rect 34257 4868 34261 4924
rect 34197 4864 34261 4868
rect 10382 4380 10446 4384
rect 10382 4324 10386 4380
rect 10386 4324 10442 4380
rect 10442 4324 10446 4380
rect 10382 4320 10446 4324
rect 10462 4380 10526 4384
rect 10462 4324 10466 4380
rect 10466 4324 10522 4380
rect 10522 4324 10526 4380
rect 10462 4320 10526 4324
rect 10542 4380 10606 4384
rect 10542 4324 10546 4380
rect 10546 4324 10602 4380
rect 10602 4324 10606 4380
rect 10542 4320 10606 4324
rect 10622 4380 10686 4384
rect 10622 4324 10626 4380
rect 10626 4324 10682 4380
rect 10682 4324 10686 4380
rect 10622 4320 10686 4324
rect 19812 4380 19876 4384
rect 19812 4324 19816 4380
rect 19816 4324 19872 4380
rect 19872 4324 19876 4380
rect 19812 4320 19876 4324
rect 19892 4380 19956 4384
rect 19892 4324 19896 4380
rect 19896 4324 19952 4380
rect 19952 4324 19956 4380
rect 19892 4320 19956 4324
rect 19972 4380 20036 4384
rect 19972 4324 19976 4380
rect 19976 4324 20032 4380
rect 20032 4324 20036 4380
rect 19972 4320 20036 4324
rect 20052 4380 20116 4384
rect 20052 4324 20056 4380
rect 20056 4324 20112 4380
rect 20112 4324 20116 4380
rect 20052 4320 20116 4324
rect 29242 4380 29306 4384
rect 29242 4324 29246 4380
rect 29246 4324 29302 4380
rect 29302 4324 29306 4380
rect 29242 4320 29306 4324
rect 29322 4380 29386 4384
rect 29322 4324 29326 4380
rect 29326 4324 29382 4380
rect 29382 4324 29386 4380
rect 29322 4320 29386 4324
rect 29402 4380 29466 4384
rect 29402 4324 29406 4380
rect 29406 4324 29462 4380
rect 29462 4324 29466 4380
rect 29402 4320 29466 4324
rect 29482 4380 29546 4384
rect 29482 4324 29486 4380
rect 29486 4324 29542 4380
rect 29542 4324 29546 4380
rect 29482 4320 29546 4324
rect 38672 4380 38736 4384
rect 38672 4324 38676 4380
rect 38676 4324 38732 4380
rect 38732 4324 38736 4380
rect 38672 4320 38736 4324
rect 38752 4380 38816 4384
rect 38752 4324 38756 4380
rect 38756 4324 38812 4380
rect 38812 4324 38816 4380
rect 38752 4320 38816 4324
rect 38832 4380 38896 4384
rect 38832 4324 38836 4380
rect 38836 4324 38892 4380
rect 38892 4324 38896 4380
rect 38832 4320 38896 4324
rect 38912 4380 38976 4384
rect 38912 4324 38916 4380
rect 38916 4324 38972 4380
rect 38972 4324 38976 4380
rect 38912 4320 38976 4324
rect 5667 3836 5731 3840
rect 5667 3780 5671 3836
rect 5671 3780 5727 3836
rect 5727 3780 5731 3836
rect 5667 3776 5731 3780
rect 5747 3836 5811 3840
rect 5747 3780 5751 3836
rect 5751 3780 5807 3836
rect 5807 3780 5811 3836
rect 5747 3776 5811 3780
rect 5827 3836 5891 3840
rect 5827 3780 5831 3836
rect 5831 3780 5887 3836
rect 5887 3780 5891 3836
rect 5827 3776 5891 3780
rect 5907 3836 5971 3840
rect 5907 3780 5911 3836
rect 5911 3780 5967 3836
rect 5967 3780 5971 3836
rect 5907 3776 5971 3780
rect 15097 3836 15161 3840
rect 15097 3780 15101 3836
rect 15101 3780 15157 3836
rect 15157 3780 15161 3836
rect 15097 3776 15161 3780
rect 15177 3836 15241 3840
rect 15177 3780 15181 3836
rect 15181 3780 15237 3836
rect 15237 3780 15241 3836
rect 15177 3776 15241 3780
rect 15257 3836 15321 3840
rect 15257 3780 15261 3836
rect 15261 3780 15317 3836
rect 15317 3780 15321 3836
rect 15257 3776 15321 3780
rect 15337 3836 15401 3840
rect 15337 3780 15341 3836
rect 15341 3780 15397 3836
rect 15397 3780 15401 3836
rect 15337 3776 15401 3780
rect 24527 3836 24591 3840
rect 24527 3780 24531 3836
rect 24531 3780 24587 3836
rect 24587 3780 24591 3836
rect 24527 3776 24591 3780
rect 24607 3836 24671 3840
rect 24607 3780 24611 3836
rect 24611 3780 24667 3836
rect 24667 3780 24671 3836
rect 24607 3776 24671 3780
rect 24687 3836 24751 3840
rect 24687 3780 24691 3836
rect 24691 3780 24747 3836
rect 24747 3780 24751 3836
rect 24687 3776 24751 3780
rect 24767 3836 24831 3840
rect 24767 3780 24771 3836
rect 24771 3780 24827 3836
rect 24827 3780 24831 3836
rect 24767 3776 24831 3780
rect 33957 3836 34021 3840
rect 33957 3780 33961 3836
rect 33961 3780 34017 3836
rect 34017 3780 34021 3836
rect 33957 3776 34021 3780
rect 34037 3836 34101 3840
rect 34037 3780 34041 3836
rect 34041 3780 34097 3836
rect 34097 3780 34101 3836
rect 34037 3776 34101 3780
rect 34117 3836 34181 3840
rect 34117 3780 34121 3836
rect 34121 3780 34177 3836
rect 34177 3780 34181 3836
rect 34117 3776 34181 3780
rect 34197 3836 34261 3840
rect 34197 3780 34201 3836
rect 34201 3780 34257 3836
rect 34257 3780 34261 3836
rect 34197 3776 34261 3780
rect 10382 3292 10446 3296
rect 10382 3236 10386 3292
rect 10386 3236 10442 3292
rect 10442 3236 10446 3292
rect 10382 3232 10446 3236
rect 10462 3292 10526 3296
rect 10462 3236 10466 3292
rect 10466 3236 10522 3292
rect 10522 3236 10526 3292
rect 10462 3232 10526 3236
rect 10542 3292 10606 3296
rect 10542 3236 10546 3292
rect 10546 3236 10602 3292
rect 10602 3236 10606 3292
rect 10542 3232 10606 3236
rect 10622 3292 10686 3296
rect 10622 3236 10626 3292
rect 10626 3236 10682 3292
rect 10682 3236 10686 3292
rect 10622 3232 10686 3236
rect 19812 3292 19876 3296
rect 19812 3236 19816 3292
rect 19816 3236 19872 3292
rect 19872 3236 19876 3292
rect 19812 3232 19876 3236
rect 19892 3292 19956 3296
rect 19892 3236 19896 3292
rect 19896 3236 19952 3292
rect 19952 3236 19956 3292
rect 19892 3232 19956 3236
rect 19972 3292 20036 3296
rect 19972 3236 19976 3292
rect 19976 3236 20032 3292
rect 20032 3236 20036 3292
rect 19972 3232 20036 3236
rect 20052 3292 20116 3296
rect 20052 3236 20056 3292
rect 20056 3236 20112 3292
rect 20112 3236 20116 3292
rect 20052 3232 20116 3236
rect 29242 3292 29306 3296
rect 29242 3236 29246 3292
rect 29246 3236 29302 3292
rect 29302 3236 29306 3292
rect 29242 3232 29306 3236
rect 29322 3292 29386 3296
rect 29322 3236 29326 3292
rect 29326 3236 29382 3292
rect 29382 3236 29386 3292
rect 29322 3232 29386 3236
rect 29402 3292 29466 3296
rect 29402 3236 29406 3292
rect 29406 3236 29462 3292
rect 29462 3236 29466 3292
rect 29402 3232 29466 3236
rect 29482 3292 29546 3296
rect 29482 3236 29486 3292
rect 29486 3236 29542 3292
rect 29542 3236 29546 3292
rect 29482 3232 29546 3236
rect 38672 3292 38736 3296
rect 38672 3236 38676 3292
rect 38676 3236 38732 3292
rect 38732 3236 38736 3292
rect 38672 3232 38736 3236
rect 38752 3292 38816 3296
rect 38752 3236 38756 3292
rect 38756 3236 38812 3292
rect 38812 3236 38816 3292
rect 38752 3232 38816 3236
rect 38832 3292 38896 3296
rect 38832 3236 38836 3292
rect 38836 3236 38892 3292
rect 38892 3236 38896 3292
rect 38832 3232 38896 3236
rect 38912 3292 38976 3296
rect 38912 3236 38916 3292
rect 38916 3236 38972 3292
rect 38972 3236 38976 3292
rect 38912 3232 38976 3236
rect 5667 2748 5731 2752
rect 5667 2692 5671 2748
rect 5671 2692 5727 2748
rect 5727 2692 5731 2748
rect 5667 2688 5731 2692
rect 5747 2748 5811 2752
rect 5747 2692 5751 2748
rect 5751 2692 5807 2748
rect 5807 2692 5811 2748
rect 5747 2688 5811 2692
rect 5827 2748 5891 2752
rect 5827 2692 5831 2748
rect 5831 2692 5887 2748
rect 5887 2692 5891 2748
rect 5827 2688 5891 2692
rect 5907 2748 5971 2752
rect 5907 2692 5911 2748
rect 5911 2692 5967 2748
rect 5967 2692 5971 2748
rect 5907 2688 5971 2692
rect 15097 2748 15161 2752
rect 15097 2692 15101 2748
rect 15101 2692 15157 2748
rect 15157 2692 15161 2748
rect 15097 2688 15161 2692
rect 15177 2748 15241 2752
rect 15177 2692 15181 2748
rect 15181 2692 15237 2748
rect 15237 2692 15241 2748
rect 15177 2688 15241 2692
rect 15257 2748 15321 2752
rect 15257 2692 15261 2748
rect 15261 2692 15317 2748
rect 15317 2692 15321 2748
rect 15257 2688 15321 2692
rect 15337 2748 15401 2752
rect 15337 2692 15341 2748
rect 15341 2692 15397 2748
rect 15397 2692 15401 2748
rect 15337 2688 15401 2692
rect 24527 2748 24591 2752
rect 24527 2692 24531 2748
rect 24531 2692 24587 2748
rect 24587 2692 24591 2748
rect 24527 2688 24591 2692
rect 24607 2748 24671 2752
rect 24607 2692 24611 2748
rect 24611 2692 24667 2748
rect 24667 2692 24671 2748
rect 24607 2688 24671 2692
rect 24687 2748 24751 2752
rect 24687 2692 24691 2748
rect 24691 2692 24747 2748
rect 24747 2692 24751 2748
rect 24687 2688 24751 2692
rect 24767 2748 24831 2752
rect 24767 2692 24771 2748
rect 24771 2692 24827 2748
rect 24827 2692 24831 2748
rect 24767 2688 24831 2692
rect 33957 2748 34021 2752
rect 33957 2692 33961 2748
rect 33961 2692 34017 2748
rect 34017 2692 34021 2748
rect 33957 2688 34021 2692
rect 34037 2748 34101 2752
rect 34037 2692 34041 2748
rect 34041 2692 34097 2748
rect 34097 2692 34101 2748
rect 34037 2688 34101 2692
rect 34117 2748 34181 2752
rect 34117 2692 34121 2748
rect 34121 2692 34177 2748
rect 34177 2692 34181 2748
rect 34117 2688 34181 2692
rect 34197 2748 34261 2752
rect 34197 2692 34201 2748
rect 34201 2692 34257 2748
rect 34257 2692 34261 2748
rect 34197 2688 34261 2692
rect 10382 2204 10446 2208
rect 10382 2148 10386 2204
rect 10386 2148 10442 2204
rect 10442 2148 10446 2204
rect 10382 2144 10446 2148
rect 10462 2204 10526 2208
rect 10462 2148 10466 2204
rect 10466 2148 10522 2204
rect 10522 2148 10526 2204
rect 10462 2144 10526 2148
rect 10542 2204 10606 2208
rect 10542 2148 10546 2204
rect 10546 2148 10602 2204
rect 10602 2148 10606 2204
rect 10542 2144 10606 2148
rect 10622 2204 10686 2208
rect 10622 2148 10626 2204
rect 10626 2148 10682 2204
rect 10682 2148 10686 2204
rect 10622 2144 10686 2148
rect 19812 2204 19876 2208
rect 19812 2148 19816 2204
rect 19816 2148 19872 2204
rect 19872 2148 19876 2204
rect 19812 2144 19876 2148
rect 19892 2204 19956 2208
rect 19892 2148 19896 2204
rect 19896 2148 19952 2204
rect 19952 2148 19956 2204
rect 19892 2144 19956 2148
rect 19972 2204 20036 2208
rect 19972 2148 19976 2204
rect 19976 2148 20032 2204
rect 20032 2148 20036 2204
rect 19972 2144 20036 2148
rect 20052 2204 20116 2208
rect 20052 2148 20056 2204
rect 20056 2148 20112 2204
rect 20112 2148 20116 2204
rect 20052 2144 20116 2148
rect 29242 2204 29306 2208
rect 29242 2148 29246 2204
rect 29246 2148 29302 2204
rect 29302 2148 29306 2204
rect 29242 2144 29306 2148
rect 29322 2204 29386 2208
rect 29322 2148 29326 2204
rect 29326 2148 29382 2204
rect 29382 2148 29386 2204
rect 29322 2144 29386 2148
rect 29402 2204 29466 2208
rect 29402 2148 29406 2204
rect 29406 2148 29462 2204
rect 29462 2148 29466 2204
rect 29402 2144 29466 2148
rect 29482 2204 29546 2208
rect 29482 2148 29486 2204
rect 29486 2148 29542 2204
rect 29542 2148 29546 2204
rect 29482 2144 29546 2148
rect 38672 2204 38736 2208
rect 38672 2148 38676 2204
rect 38676 2148 38732 2204
rect 38732 2148 38736 2204
rect 38672 2144 38736 2148
rect 38752 2204 38816 2208
rect 38752 2148 38756 2204
rect 38756 2148 38812 2204
rect 38812 2148 38816 2204
rect 38752 2144 38816 2148
rect 38832 2204 38896 2208
rect 38832 2148 38836 2204
rect 38836 2148 38892 2204
rect 38892 2148 38896 2204
rect 38832 2144 38896 2148
rect 38912 2204 38976 2208
rect 38912 2148 38916 2204
rect 38916 2148 38972 2204
rect 38972 2148 38976 2204
rect 38912 2144 38976 2148
<< metal4 >>
rect 5659 9280 5979 9840
rect 5659 9216 5667 9280
rect 5731 9216 5747 9280
rect 5811 9216 5827 9280
rect 5891 9216 5907 9280
rect 5971 9216 5979 9280
rect 5659 8192 5979 9216
rect 5659 8128 5667 8192
rect 5731 8128 5747 8192
rect 5811 8128 5827 8192
rect 5891 8128 5907 8192
rect 5971 8128 5979 8192
rect 5659 7104 5979 8128
rect 5659 7040 5667 7104
rect 5731 7040 5747 7104
rect 5811 7040 5827 7104
rect 5891 7040 5907 7104
rect 5971 7040 5979 7104
rect 5659 6016 5979 7040
rect 5659 5952 5667 6016
rect 5731 5952 5747 6016
rect 5811 5952 5827 6016
rect 5891 5952 5907 6016
rect 5971 5952 5979 6016
rect 5659 4928 5979 5952
rect 5659 4864 5667 4928
rect 5731 4864 5747 4928
rect 5811 4864 5827 4928
rect 5891 4864 5907 4928
rect 5971 4864 5979 4928
rect 5659 3840 5979 4864
rect 5659 3776 5667 3840
rect 5731 3776 5747 3840
rect 5811 3776 5827 3840
rect 5891 3776 5907 3840
rect 5971 3776 5979 3840
rect 5659 2752 5979 3776
rect 5659 2688 5667 2752
rect 5731 2688 5747 2752
rect 5811 2688 5827 2752
rect 5891 2688 5907 2752
rect 5971 2688 5979 2752
rect 5659 2128 5979 2688
rect 10374 9824 10694 9840
rect 10374 9760 10382 9824
rect 10446 9760 10462 9824
rect 10526 9760 10542 9824
rect 10606 9760 10622 9824
rect 10686 9760 10694 9824
rect 10374 8736 10694 9760
rect 10374 8672 10382 8736
rect 10446 8672 10462 8736
rect 10526 8672 10542 8736
rect 10606 8672 10622 8736
rect 10686 8672 10694 8736
rect 10374 7648 10694 8672
rect 10374 7584 10382 7648
rect 10446 7584 10462 7648
rect 10526 7584 10542 7648
rect 10606 7584 10622 7648
rect 10686 7584 10694 7648
rect 10374 6560 10694 7584
rect 10374 6496 10382 6560
rect 10446 6496 10462 6560
rect 10526 6496 10542 6560
rect 10606 6496 10622 6560
rect 10686 6496 10694 6560
rect 10374 5472 10694 6496
rect 10374 5408 10382 5472
rect 10446 5408 10462 5472
rect 10526 5408 10542 5472
rect 10606 5408 10622 5472
rect 10686 5408 10694 5472
rect 10374 4384 10694 5408
rect 10374 4320 10382 4384
rect 10446 4320 10462 4384
rect 10526 4320 10542 4384
rect 10606 4320 10622 4384
rect 10686 4320 10694 4384
rect 10374 3296 10694 4320
rect 10374 3232 10382 3296
rect 10446 3232 10462 3296
rect 10526 3232 10542 3296
rect 10606 3232 10622 3296
rect 10686 3232 10694 3296
rect 10374 2208 10694 3232
rect 10374 2144 10382 2208
rect 10446 2144 10462 2208
rect 10526 2144 10542 2208
rect 10606 2144 10622 2208
rect 10686 2144 10694 2208
rect 10374 2128 10694 2144
rect 15089 9280 15409 9840
rect 15089 9216 15097 9280
rect 15161 9216 15177 9280
rect 15241 9216 15257 9280
rect 15321 9216 15337 9280
rect 15401 9216 15409 9280
rect 15089 8192 15409 9216
rect 15089 8128 15097 8192
rect 15161 8128 15177 8192
rect 15241 8128 15257 8192
rect 15321 8128 15337 8192
rect 15401 8128 15409 8192
rect 15089 7104 15409 8128
rect 15089 7040 15097 7104
rect 15161 7040 15177 7104
rect 15241 7040 15257 7104
rect 15321 7040 15337 7104
rect 15401 7040 15409 7104
rect 15089 6016 15409 7040
rect 15089 5952 15097 6016
rect 15161 5952 15177 6016
rect 15241 5952 15257 6016
rect 15321 5952 15337 6016
rect 15401 5952 15409 6016
rect 15089 4928 15409 5952
rect 15089 4864 15097 4928
rect 15161 4864 15177 4928
rect 15241 4864 15257 4928
rect 15321 4864 15337 4928
rect 15401 4864 15409 4928
rect 15089 3840 15409 4864
rect 15089 3776 15097 3840
rect 15161 3776 15177 3840
rect 15241 3776 15257 3840
rect 15321 3776 15337 3840
rect 15401 3776 15409 3840
rect 15089 2752 15409 3776
rect 15089 2688 15097 2752
rect 15161 2688 15177 2752
rect 15241 2688 15257 2752
rect 15321 2688 15337 2752
rect 15401 2688 15409 2752
rect 15089 2128 15409 2688
rect 19804 9824 20124 9840
rect 19804 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20052 9824
rect 20116 9760 20124 9824
rect 19804 8736 20124 9760
rect 19804 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20052 8736
rect 20116 8672 20124 8736
rect 19804 7648 20124 8672
rect 19804 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20052 7648
rect 20116 7584 20124 7648
rect 19804 6560 20124 7584
rect 19804 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20052 6560
rect 20116 6496 20124 6560
rect 19804 5472 20124 6496
rect 19804 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20052 5472
rect 20116 5408 20124 5472
rect 19804 4384 20124 5408
rect 19804 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20052 4384
rect 20116 4320 20124 4384
rect 19804 3296 20124 4320
rect 19804 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20052 3296
rect 20116 3232 20124 3296
rect 19804 2208 20124 3232
rect 19804 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20052 2208
rect 20116 2144 20124 2208
rect 19804 2128 20124 2144
rect 24519 9280 24839 9840
rect 24519 9216 24527 9280
rect 24591 9216 24607 9280
rect 24671 9216 24687 9280
rect 24751 9216 24767 9280
rect 24831 9216 24839 9280
rect 24519 8192 24839 9216
rect 24519 8128 24527 8192
rect 24591 8128 24607 8192
rect 24671 8128 24687 8192
rect 24751 8128 24767 8192
rect 24831 8128 24839 8192
rect 24519 7104 24839 8128
rect 24519 7040 24527 7104
rect 24591 7040 24607 7104
rect 24671 7040 24687 7104
rect 24751 7040 24767 7104
rect 24831 7040 24839 7104
rect 24519 6016 24839 7040
rect 24519 5952 24527 6016
rect 24591 5952 24607 6016
rect 24671 5952 24687 6016
rect 24751 5952 24767 6016
rect 24831 5952 24839 6016
rect 24519 4928 24839 5952
rect 24519 4864 24527 4928
rect 24591 4864 24607 4928
rect 24671 4864 24687 4928
rect 24751 4864 24767 4928
rect 24831 4864 24839 4928
rect 24519 3840 24839 4864
rect 24519 3776 24527 3840
rect 24591 3776 24607 3840
rect 24671 3776 24687 3840
rect 24751 3776 24767 3840
rect 24831 3776 24839 3840
rect 24519 2752 24839 3776
rect 24519 2688 24527 2752
rect 24591 2688 24607 2752
rect 24671 2688 24687 2752
rect 24751 2688 24767 2752
rect 24831 2688 24839 2752
rect 24519 2128 24839 2688
rect 29234 9824 29554 9840
rect 29234 9760 29242 9824
rect 29306 9760 29322 9824
rect 29386 9760 29402 9824
rect 29466 9760 29482 9824
rect 29546 9760 29554 9824
rect 29234 8736 29554 9760
rect 29234 8672 29242 8736
rect 29306 8672 29322 8736
rect 29386 8672 29402 8736
rect 29466 8672 29482 8736
rect 29546 8672 29554 8736
rect 29234 7648 29554 8672
rect 29234 7584 29242 7648
rect 29306 7584 29322 7648
rect 29386 7584 29402 7648
rect 29466 7584 29482 7648
rect 29546 7584 29554 7648
rect 29234 6560 29554 7584
rect 29234 6496 29242 6560
rect 29306 6496 29322 6560
rect 29386 6496 29402 6560
rect 29466 6496 29482 6560
rect 29546 6496 29554 6560
rect 29234 5472 29554 6496
rect 29234 5408 29242 5472
rect 29306 5408 29322 5472
rect 29386 5408 29402 5472
rect 29466 5408 29482 5472
rect 29546 5408 29554 5472
rect 29234 4384 29554 5408
rect 29234 4320 29242 4384
rect 29306 4320 29322 4384
rect 29386 4320 29402 4384
rect 29466 4320 29482 4384
rect 29546 4320 29554 4384
rect 29234 3296 29554 4320
rect 29234 3232 29242 3296
rect 29306 3232 29322 3296
rect 29386 3232 29402 3296
rect 29466 3232 29482 3296
rect 29546 3232 29554 3296
rect 29234 2208 29554 3232
rect 29234 2144 29242 2208
rect 29306 2144 29322 2208
rect 29386 2144 29402 2208
rect 29466 2144 29482 2208
rect 29546 2144 29554 2208
rect 29234 2128 29554 2144
rect 33949 9280 34269 9840
rect 33949 9216 33957 9280
rect 34021 9216 34037 9280
rect 34101 9216 34117 9280
rect 34181 9216 34197 9280
rect 34261 9216 34269 9280
rect 33949 8192 34269 9216
rect 33949 8128 33957 8192
rect 34021 8128 34037 8192
rect 34101 8128 34117 8192
rect 34181 8128 34197 8192
rect 34261 8128 34269 8192
rect 33949 7104 34269 8128
rect 33949 7040 33957 7104
rect 34021 7040 34037 7104
rect 34101 7040 34117 7104
rect 34181 7040 34197 7104
rect 34261 7040 34269 7104
rect 33949 6016 34269 7040
rect 33949 5952 33957 6016
rect 34021 5952 34037 6016
rect 34101 5952 34117 6016
rect 34181 5952 34197 6016
rect 34261 5952 34269 6016
rect 33949 4928 34269 5952
rect 33949 4864 33957 4928
rect 34021 4864 34037 4928
rect 34101 4864 34117 4928
rect 34181 4864 34197 4928
rect 34261 4864 34269 4928
rect 33949 3840 34269 4864
rect 33949 3776 33957 3840
rect 34021 3776 34037 3840
rect 34101 3776 34117 3840
rect 34181 3776 34197 3840
rect 34261 3776 34269 3840
rect 33949 2752 34269 3776
rect 33949 2688 33957 2752
rect 34021 2688 34037 2752
rect 34101 2688 34117 2752
rect 34181 2688 34197 2752
rect 34261 2688 34269 2752
rect 33949 2128 34269 2688
rect 38664 9824 38984 9840
rect 38664 9760 38672 9824
rect 38736 9760 38752 9824
rect 38816 9760 38832 9824
rect 38896 9760 38912 9824
rect 38976 9760 38984 9824
rect 38664 8736 38984 9760
rect 38664 8672 38672 8736
rect 38736 8672 38752 8736
rect 38816 8672 38832 8736
rect 38896 8672 38912 8736
rect 38976 8672 38984 8736
rect 38664 7648 38984 8672
rect 38664 7584 38672 7648
rect 38736 7584 38752 7648
rect 38816 7584 38832 7648
rect 38896 7584 38912 7648
rect 38976 7584 38984 7648
rect 38664 6560 38984 7584
rect 38664 6496 38672 6560
rect 38736 6496 38752 6560
rect 38816 6496 38832 6560
rect 38896 6496 38912 6560
rect 38976 6496 38984 6560
rect 38664 5472 38984 6496
rect 38664 5408 38672 5472
rect 38736 5408 38752 5472
rect 38816 5408 38832 5472
rect 38896 5408 38912 5472
rect 38976 5408 38984 5472
rect 38664 4384 38984 5408
rect 38664 4320 38672 4384
rect 38736 4320 38752 4384
rect 38816 4320 38832 4384
rect 38896 4320 38912 4384
rect 38976 4320 38984 4384
rect 38664 3296 38984 4320
rect 38664 3232 38672 3296
rect 38736 3232 38752 3296
rect 38816 3232 38832 3296
rect 38896 3232 38912 3296
rect 38976 3232 38984 3296
rect 38664 2208 38984 3232
rect 38664 2144 38672 2208
rect 38736 2144 38752 2208
rect 38816 2144 38832 2208
rect 38896 2144 38912 2208
rect 38976 2144 38984 2208
rect 38664 2128 38984 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_20
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_286
timestamp 1688980957
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_298
timestamp 1688980957
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_306
timestamp 1688980957
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_314
timestamp 1688980957
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_326
timestamp 1688980957
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_334
timestamp 1688980957
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_342
timestamp 1688980957
transform 1 0 32568 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_354
timestamp 1688980957
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_362
timestamp 1688980957
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_370
timestamp 1688980957
transform 1 0 35144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_382
timestamp 1688980957
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1688980957
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_398 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37720 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_6
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_18
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_30
timestamp 1688980957
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_42
timestamp 1688980957
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1688980957
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1688980957
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_401
timestamp 1688980957
transform 1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1688980957
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_6
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_13
timestamp 1688980957
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_25
timestamp 1688980957
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_153
timestamp 1688980957
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_160
timestamp 1688980957
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_188
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_209
timestamp 1688980957
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_216
timestamp 1688980957
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_244
timestamp 1688980957
transform 1 0 23552 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_265
timestamp 1688980957
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_307
timestamp 1688980957
transform 1 0 29348 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_321
timestamp 1688980957
transform 1 0 30636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_357
timestamp 1688980957
transform 1 0 33948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_363
timestamp 1688980957
transform 1 0 34500 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_365
timestamp 1688980957
transform 1 0 34684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_377
timestamp 1688980957
transform 1 0 35788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_401
timestamp 1688980957
transform 1 0 37996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_2
timestamp 1688980957
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_3
timestamp 1688980957
transform -1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_4
timestamp 1688980957
transform -1 0 29348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_5
timestamp 1688980957
transform -1 0 31924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_6
timestamp 1688980957
transform -1 0 18400 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_7
timestamp 1688980957
transform -1 0 24196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_8
timestamp 1688980957
transform -1 0 21620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_9
timestamp 1688980957
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_10
timestamp 1688980957
transform 1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_11
timestamp 1688980957
transform -1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_12
timestamp 1688980957
transform -1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_13
timestamp 1688980957
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_14
timestamp 1688980957
transform 1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_15
timestamp 1688980957
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_16
timestamp 1688980957
transform -1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_17
timestamp 1688980957
transform -1 0 19044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_18
timestamp 1688980957
transform 1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_19
timestamp 1688980957
transform -1 0 23552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_20
timestamp 1688980957
transform -1 0 26128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_21
timestamp 1688980957
transform -1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_22
timestamp 1688980957
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_23
timestamp 1688980957
transform -1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_24
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_25
timestamp 1688980957
transform -1 0 38548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_26
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_27
timestamp 1688980957
transform 1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_28
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_29
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_30
timestamp 1688980957
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_31
timestamp 1688980957
transform 1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_32
timestamp 1688980957
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_33
timestamp 1688980957
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_34
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_35
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_36
timestamp 1688980957
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_37
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ioenb_38
timestamp 1688980957
transform -1 0 38548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 0 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_oeb[10]
port 1 nsew signal tristate
flabel metal2 s 7102 11200 7158 12000 0 FreeSans 224 90 0 0 io_oeb[11]
port 2 nsew signal tristate
flabel metal2 s 34150 11200 34206 12000 0 FreeSans 224 90 0 0 io_oeb[12]
port 3 nsew signal tristate
flabel metal2 s 28998 11200 29054 12000 0 FreeSans 224 90 0 0 io_oeb[13]
port 4 nsew signal tristate
flabel metal2 s 31574 11200 31630 12000 0 FreeSans 224 90 0 0 io_oeb[14]
port 5 nsew signal tristate
flabel metal2 s 18050 11200 18106 12000 0 FreeSans 224 90 0 0 io_oeb[15]
port 6 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 7 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 8 nsew signal tristate
flabel metal2 s 4526 11200 4582 12000 0 FreeSans 224 90 0 0 io_oeb[18]
port 9 nsew signal tristate
flabel metal3 s 39200 3408 40000 3528 0 FreeSans 480 0 0 0 io_oeb[19]
port 10 nsew signal tristate
flabel metal2 s 20626 11200 20682 12000 0 FreeSans 224 90 0 0 io_oeb[1]
port 11 nsew signal tristate
flabel metal2 s 9678 11200 9734 12000 0 FreeSans 224 90 0 0 io_oeb[20]
port 12 nsew signal tristate
flabel metal2 s 1950 11200 2006 12000 0 FreeSans 224 90 0 0 io_oeb[21]
port 13 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 14 nsew signal tristate
flabel metal3 s 39200 688 40000 808 0 FreeSans 480 0 0 0 io_oeb[23]
port 15 nsew signal tristate
flabel metal3 s 39200 6128 40000 6248 0 FreeSans 480 0 0 0 io_oeb[24]
port 16 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 17 nsew signal tristate
flabel metal2 s 15474 11200 15530 12000 0 FreeSans 224 90 0 0 io_oeb[26]
port 18 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 io_oeb[27]
port 19 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 20 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 21 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 22 nsew signal tristate
flabel metal2 s 36726 11200 36782 12000 0 FreeSans 224 90 0 0 io_oeb[30]
port 23 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 24 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 25 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 26 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 io_oeb[34]
port 27 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 28 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 29 nsew signal tristate
flabel metal3 s 39200 8848 40000 8968 0 FreeSans 480 0 0 0 io_oeb[37]
port 30 nsew signal tristate
flabel metal2 s 39302 11200 39358 12000 0 FreeSans 224 90 0 0 io_oeb[3]
port 31 nsew signal tristate
flabel metal2 s 23202 11200 23258 12000 0 FreeSans 224 90 0 0 io_oeb[4]
port 32 nsew signal tristate
flabel metal2 s 25778 11200 25834 12000 0 FreeSans 224 90 0 0 io_oeb[5]
port 33 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 34 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_oeb[7]
port 35 nsew signal tristate
flabel metal2 s 12254 11200 12310 12000 0 FreeSans 224 90 0 0 io_oeb[8]
port 36 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 37 nsew signal tristate
flabel metal4 s 5659 2128 5979 9840 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 15089 2128 15409 9840 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 24519 2128 24839 9840 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 33949 2128 34269 9840 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 10374 2128 10694 9840 0 FreeSans 1920 90 0 0 vssd1
port 39 nsew ground bidirectional
flabel metal4 s 19804 2128 20124 9840 0 FreeSans 1920 90 0 0 vssd1
port 39 nsew ground bidirectional
flabel metal4 s 29234 2128 29554 9840 0 FreeSans 1920 90 0 0 vssd1
port 39 nsew ground bidirectional
flabel metal4 s 38664 2128 38984 9840 0 FreeSans 1920 90 0 0 vssd1
port 39 nsew ground bidirectional
rlabel metal1 19964 9248 19964 9248 0 vccd1
rlabel via1 20044 9792 20044 9792 0 vssd1
rlabel metal2 37398 1027 37398 1027 0 net1
rlabel via2 38502 3485 38502 3485 0 net10
rlabel metal2 9798 9607 9798 9607 0 net11
rlabel metal2 2070 9607 2070 9607 0 net12
rlabel metal2 27094 1027 27094 1027 0 net13
rlabel metal2 38502 1581 38502 1581 0 net14
rlabel metal2 13570 1027 13570 1027 0 net15
rlabel metal2 20700 9660 20700 9660 0 net16
rlabel metal2 18722 1027 18722 1027 0 net17
rlabel metal2 38870 11220 38870 11220 0 net18
rlabel metal2 23322 9607 23322 9607 0 net19
rlabel metal3 1050 8228 1050 8228 0 net2
rlabel metal2 25898 9607 25898 9607 0 net20
rlabel metal2 16146 1027 16146 1027 0 net21
rlabel metal1 2116 9486 2116 9486 0 net22
rlabel metal2 12374 9607 12374 9607 0 net23
rlabel via1 34270 9641 34270 9641 0 net24
rlabel via2 38502 6205 38502 6205 0 net25
rlabel metal2 46 823 46 823 0 net26
rlabel via1 15594 9641 15594 9641 0 net27
rlabel metal3 820 2788 820 2788 0 net28
rlabel metal2 7774 959 7774 959 0 net29
rlabel metal2 7222 9607 7222 9607 0 net3
rlabel metal2 34822 959 34822 959 0 net30
rlabel via1 36846 9641 36846 9641 0 net31
rlabel metal2 29670 959 29670 959 0 net32
rlabel metal2 2622 959 2622 959 0 net33
rlabel metal2 5198 959 5198 959 0 net34
rlabel metal3 1050 5508 1050 5508 0 net35
rlabel metal2 32246 959 32246 959 0 net36
rlabel metal2 10350 823 10350 823 0 net37
rlabel via2 38502 8891 38502 8891 0 net38
rlabel metal2 29118 9607 29118 9607 0 net4
rlabel metal2 31694 9607 31694 9607 0 net5
rlabel metal2 18170 9607 18170 9607 0 net6
rlabel metal2 23874 1027 23874 1027 0 net7
rlabel metal2 21298 1027 21298 1027 0 net8
rlabel metal2 4646 9607 4646 9607 0 net9
<< properties >>
string FIXED_BBOX 0 0 40000 12000
<< end >>
