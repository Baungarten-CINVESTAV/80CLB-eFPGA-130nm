// This is the unpowered netlist.
module sb_1__1_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
    ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
 input [8:0] chanx_left_in;
 output [8:0] chanx_left_out;
 input [8:0] chanx_right_in;
 output [8:0] chanx_right_out;
 input [8:0] chany_bottom_in;
 output [8:0] chany_bottom_out;
 input [8:0] chany_top_in;
 output [8:0] chany_top_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire clknet_0_prog_clk;
 wire clknet_2_0__leaf_prog_clk;
 wire clknet_2_1__leaf_prog_clk;
 wire clknet_2_2__leaf_prog_clk;
 wire clknet_2_3__leaf_prog_clk;
 wire \mem_bottom_track_1.DFF_0_.D ;
 wire \mem_bottom_track_1.DFF_0_.Q ;
 wire \mem_bottom_track_1.DFF_1_.Q ;
 wire \mem_bottom_track_1.DFF_2_.Q ;
 wire \mem_bottom_track_1.DFF_3_.Q ;
 wire \mem_bottom_track_17.DFF_0_.D ;
 wire \mem_bottom_track_17.DFF_0_.Q ;
 wire \mem_bottom_track_17.DFF_1_.Q ;
 wire \mem_bottom_track_17.DFF_2_.Q ;
 wire \mem_bottom_track_17.DFF_3_.Q ;
 wire \mem_bottom_track_9.DFF_0_.Q ;
 wire \mem_bottom_track_9.DFF_1_.Q ;
 wire \mem_bottom_track_9.DFF_2_.Q ;
 wire \mem_left_track_1.DFF_0_.Q ;
 wire \mem_left_track_1.DFF_1_.Q ;
 wire \mem_left_track_1.DFF_2_.Q ;
 wire \mem_left_track_1.DFF_3_.Q ;
 wire \mem_left_track_17.DFF_0_.D ;
 wire \mem_left_track_17.DFF_0_.Q ;
 wire \mem_left_track_17.DFF_1_.Q ;
 wire \mem_left_track_17.DFF_2_.Q ;
 wire \mem_left_track_9.DFF_0_.Q ;
 wire \mem_left_track_9.DFF_1_.Q ;
 wire \mem_left_track_9.DFF_2_.Q ;
 wire \mem_right_track_0.DFF_0_.D ;
 wire \mem_right_track_0.DFF_0_.Q ;
 wire \mem_right_track_0.DFF_1_.Q ;
 wire \mem_right_track_0.DFF_2_.Q ;
 wire \mem_right_track_0.DFF_3_.Q ;
 wire \mem_right_track_16.DFF_0_.D ;
 wire \mem_right_track_16.DFF_0_.Q ;
 wire \mem_right_track_16.DFF_1_.Q ;
 wire \mem_right_track_16.DFF_2_.Q ;
 wire \mem_right_track_8.DFF_0_.Q ;
 wire \mem_right_track_8.DFF_1_.Q ;
 wire \mem_right_track_8.DFF_2_.Q ;
 wire \mem_top_track_0.DFF_0_.Q ;
 wire \mem_top_track_0.DFF_1_.Q ;
 wire \mem_top_track_0.DFF_2_.Q ;
 wire \mem_top_track_0.DFF_3_.Q ;
 wire \mem_top_track_16.DFF_0_.D ;
 wire \mem_top_track_16.DFF_0_.Q ;
 wire \mem_top_track_16.DFF_1_.Q ;
 wire \mem_top_track_16.DFF_2_.Q ;
 wire \mem_top_track_8.DFF_0_.Q ;
 wire \mem_top_track_8.DFF_1_.Q ;
 wire \mem_top_track_8.DFF_2_.Q ;
 wire \mux_bottom_track_1.INVTX1_0_.out ;
 wire \mux_bottom_track_1.INVTX1_1_.out ;
 wire \mux_bottom_track_1.INVTX1_2_.out ;
 wire \mux_bottom_track_1.INVTX1_3_.out ;
 wire \mux_bottom_track_1.INVTX1_4_.out ;
 wire \mux_bottom_track_1.INVTX1_5_.out ;
 wire \mux_bottom_track_1.INVTX1_6_.out ;
 wire \mux_bottom_track_1.INVTX1_7_.out ;
 wire \mux_bottom_track_1.INVTX1_8_.out ;
 wire \mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_1.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_17.INVTX1_0_.out ;
 wire \mux_bottom_track_17.INVTX1_1_.out ;
 wire \mux_bottom_track_17.INVTX1_2_.out ;
 wire \mux_bottom_track_17.INVTX1_3_.out ;
 wire \mux_bottom_track_17.INVTX1_4_.out ;
 wire \mux_bottom_track_17.INVTX1_5_.out ;
 wire \mux_bottom_track_17.INVTX1_6_.out ;
 wire \mux_bottom_track_17.INVTX1_7_.out ;
 wire \mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_17.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_9.INVTX1_0_.out ;
 wire \mux_bottom_track_9.INVTX1_1_.out ;
 wire \mux_bottom_track_9.INVTX1_2_.out ;
 wire \mux_bottom_track_9.INVTX1_3_.out ;
 wire \mux_bottom_track_9.INVTX1_4_.out ;
 wire \mux_bottom_track_9.INVTX1_5_.out ;
 wire \mux_bottom_track_9.INVTX1_6_.out ;
 wire \mux_bottom_track_9.INVTX1_7_.out ;
 wire \mux_bottom_track_9.INVTX1_8_.out ;
 wire \mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_bottom_track_9.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_left_track_1.INVTX1_1_.out ;
 wire \mux_left_track_1.INVTX1_5_.out ;
 wire \mux_left_track_1.INVTX1_6_.out ;
 wire \mux_left_track_1.INVTX1_7_.out ;
 wire \mux_left_track_1.INVTX1_8_.out ;
 wire \mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_left_track_1.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_left_track_17.INVTX1_2_.out ;
 wire \mux_left_track_17.INVTX1_5_.out ;
 wire \mux_left_track_17.INVTX1_6_.out ;
 wire \mux_left_track_17.INVTX1_7_.out ;
 wire \mux_left_track_17.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_left_track_17.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_left_track_9.INVTX1_2_.out ;
 wire \mux_left_track_9.INVTX1_5_.out ;
 wire \mux_left_track_9.INVTX1_6_.out ;
 wire \mux_left_track_9.INVTX1_7_.out ;
 wire \mux_left_track_9.INVTX1_8_.out ;
 wire \mux_left_track_9.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_left_track_9.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_right_track_0.INVTX1_3_.out ;
 wire \mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_right_track_0.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_right_track_16.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_right_track_8.INVTX1_3_.out ;
 wire \mux_right_track_8.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_right_track_8.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_top_track_0.INVTX1_0_.out ;
 wire \mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_top_track_0.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_top_track_16.mux_l4_in_0_.TGATE_0_.out ;
 wire \mux_top_track_8.INVTX1_0_.out ;
 wire \mux_top_track_8.mux_l1_in_0_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l1_in_1_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l2_in_0_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l2_in_1_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l2_in_2_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l2_in_3_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l3_in_0_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l3_in_1_.TGATE_0_.out ;
 wire \mux_top_track_8.mux_l4_in_0_.TGATE_0_.out ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__fill_1 FILLER_0_0_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__clkbuf_1 _324_ (.A(\mem_bottom_track_1.DFF_0_.Q ),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _325_ (.A(_060_),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _326_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _327_ (.A(_061_),
    .X(_182_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(\mem_bottom_track_1.DFF_0_.Q ),
    .Y(_192_));
 sky130_fd_sc_hd__clkbuf_1 _329_ (.A(\mem_bottom_track_1.DFF_0_.Q ),
    .X(_062_));
 sky130_fd_sc_hd__clkbuf_1 _330_ (.A(_062_),
    .X(_183_));
 sky130_fd_sc_hd__clkbuf_1 _331_ (.A(\mem_bottom_track_1.DFF_2_.Q ),
    .X(_063_));
 sky130_fd_sc_hd__clkbuf_1 _332_ (.A(_063_),
    .X(_178_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .Y(_190_));
 sky130_fd_sc_hd__clkbuf_1 _334_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .X(_064_));
 sky130_fd_sc_hd__clkbuf_1 _335_ (.A(_064_),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_1 _336_ (.A(\mem_bottom_track_1.DFF_3_.Q ),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_1 _337_ (.A(_065_),
    .X(_176_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\mem_bottom_track_1.DFF_2_.Q ),
    .Y(_186_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .Y(_189_));
 sky130_fd_sc_hd__clkbuf_1 _340_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .X(_066_));
 sky130_fd_sc_hd__clkbuf_1 _341_ (.A(_066_),
    .X(_180_));
 sky130_fd_sc_hd__clkbuf_1 _342_ (.A(\mem_bottom_track_1.DFF_2_.Q ),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_1 _343_ (.A(_067_),
    .X(_177_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .Y(_188_));
 sky130_fd_sc_hd__clkbuf_1 _345_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .X(_068_));
 sky130_fd_sc_hd__clkbuf_1 _346_ (.A(_068_),
    .X(_179_));
 sky130_fd_sc_hd__inv_2 _347_ (.A(\mem_right_track_16.DFF_0_.D ),
    .Y(_167_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(\mem_right_track_8.DFF_2_.Q ),
    .Y(_169_));
 sky130_fd_sc_hd__inv_2 _349_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .Y(_173_));
 sky130_fd_sc_hd__inv_2 _350_ (.A(\mem_right_track_8.DFF_0_.Q ),
    .Y(_175_));
 sky130_fd_sc_hd__clkbuf_1 _351_ (.A(\mem_right_track_8.DFF_0_.Q ),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _352_ (.A(_069_),
    .X(_166_));
 sky130_fd_sc_hd__clkbuf_1 _353_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _354_ (.A(_070_),
    .X(_164_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(\mem_right_track_8.DFF_0_.Q ),
    .Y(_174_));
 sky130_fd_sc_hd__clkbuf_1 _356_ (.A(\mem_right_track_8.DFF_0_.Q ),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _357_ (.A(_071_),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_1 _358_ (.A(\mem_right_track_8.DFF_2_.Q ),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_1 _359_ (.A(_072_),
    .X(_160_));
 sky130_fd_sc_hd__inv_2 _360_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .Y(_172_));
 sky130_fd_sc_hd__clkbuf_1 _361_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(_073_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _363_ (.A(\mem_right_track_16.DFF_0_.D ),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _364_ (.A(_074_),
    .X(_158_));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\mem_right_track_8.DFF_2_.Q ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_2 _366_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .Y(_171_));
 sky130_fd_sc_hd__clkbuf_1 _367_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _368_ (.A(_075_),
    .X(_162_));
 sky130_fd_sc_hd__clkbuf_1 _369_ (.A(\mem_right_track_8.DFF_2_.Q ),
    .X(_076_));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(_076_),
    .X(_159_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .Y(_170_));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(\mem_right_track_8.DFF_1_.Q ),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_1 _373_ (.A(_077_),
    .X(_161_));
 sky130_fd_sc_hd__inv_2 _374_ (.A(\mem_right_track_0.DFF_3_.Q ),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(\mem_right_track_0.DFF_2_.Q ),
    .Y(_151_));
 sky130_fd_sc_hd__inv_2 _376_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(\mem_right_track_0.DFF_0_.Q ),
    .Y(_157_));
 sky130_fd_sc_hd__clkbuf_1 _378_ (.A(\mem_right_track_0.DFF_0_.Q ),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_078_),
    .X(_148_));
 sky130_fd_sc_hd__clkbuf_1 _380_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .X(_079_));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(_079_),
    .X(_146_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(\mem_right_track_0.DFF_0_.Q ),
    .Y(_156_));
 sky130_fd_sc_hd__clkbuf_1 _383_ (.A(\mem_right_track_0.DFF_0_.Q ),
    .X(_080_));
 sky130_fd_sc_hd__clkbuf_1 _384_ (.A(_080_),
    .X(_147_));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(\mem_right_track_0.DFF_2_.Q ),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_1 _386_ (.A(_081_),
    .X(_142_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .Y(_154_));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .X(_082_));
 sky130_fd_sc_hd__clkbuf_1 _389_ (.A(_082_),
    .X(_145_));
 sky130_fd_sc_hd__clkbuf_1 _390_ (.A(\mem_right_track_0.DFF_3_.Q ),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_1 _391_ (.A(_083_),
    .X(_140_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(\mem_right_track_0.DFF_2_.Q ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .Y(_153_));
 sky130_fd_sc_hd__clkbuf_1 _394_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_1 _395_ (.A(_084_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(\mem_right_track_0.DFF_2_.Q ),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_1 _397_ (.A(_085_),
    .X(_141_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .Y(_152_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(\mem_right_track_0.DFF_1_.Q ),
    .X(_086_));
 sky130_fd_sc_hd__clkbuf_1 _400_ (.A(_086_),
    .X(_143_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(\mem_top_track_16.DFF_0_.D ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(\mem_top_track_8.DFF_2_.Q ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _403_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(\mem_top_track_8.DFF_0_.Q ),
    .Y(_139_));
 sky130_fd_sc_hd__clkbuf_1 _405_ (.A(\mem_top_track_8.DFF_0_.Q ),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_1 _406_ (.A(_087_),
    .X(_130_));
 sky130_fd_sc_hd__clkbuf_1 _407_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .X(_088_));
 sky130_fd_sc_hd__clkbuf_1 _408_ (.A(_088_),
    .X(_128_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(\mem_top_track_8.DFF_0_.Q ),
    .Y(_138_));
 sky130_fd_sc_hd__clkbuf_1 _410_ (.A(\mem_top_track_8.DFF_0_.Q ),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_1 _411_ (.A(_089_),
    .X(_129_));
 sky130_fd_sc_hd__clkbuf_1 _412_ (.A(\mem_top_track_8.DFF_2_.Q ),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _413_ (.A(_090_),
    .X(_124_));
 sky130_fd_sc_hd__inv_2 _414_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .Y(_136_));
 sky130_fd_sc_hd__clkbuf_1 _415_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .X(_091_));
 sky130_fd_sc_hd__clkbuf_1 _416_ (.A(_091_),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _417_ (.A(\mem_top_track_16.DFF_0_.D ),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_1 _418_ (.A(_092_),
    .X(_122_));
 sky130_fd_sc_hd__inv_2 _419_ (.A(\mem_top_track_8.DFF_2_.Q ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .Y(_135_));
 sky130_fd_sc_hd__clkbuf_1 _421_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .X(_093_));
 sky130_fd_sc_hd__clkbuf_1 _422_ (.A(_093_),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _423_ (.A(\mem_top_track_8.DFF_2_.Q ),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_094_),
    .X(_123_));
 sky130_fd_sc_hd__inv_2 _425_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .Y(_134_));
 sky130_fd_sc_hd__clkbuf_1 _426_ (.A(\mem_top_track_8.DFF_1_.Q ),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_1 _427_ (.A(_095_),
    .X(_125_));
 sky130_fd_sc_hd__inv_2 _428_ (.A(\mem_top_track_0.DFF_2_.Q ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(\mem_top_track_0.DFF_3_.Q ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(\mem_top_track_0.DFF_2_.Q ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(\mem_top_track_0.DFF_0_.Q ),
    .Y(_121_));
 sky130_fd_sc_hd__clkbuf_1 _434_ (.A(\mem_top_track_0.DFF_0_.Q ),
    .X(_096_));
 sky130_fd_sc_hd__clkbuf_1 _435_ (.A(_096_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _436_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .X(_097_));
 sky130_fd_sc_hd__clkbuf_1 _437_ (.A(_097_),
    .X(_110_));
 sky130_fd_sc_hd__inv_2 _438_ (.A(\mem_top_track_0.DFF_0_.Q ),
    .Y(_120_));
 sky130_fd_sc_hd__clkbuf_1 _439_ (.A(\mem_top_track_0.DFF_0_.Q ),
    .X(_098_));
 sky130_fd_sc_hd__clkbuf_1 _440_ (.A(_098_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _441_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .X(_099_));
 sky130_fd_sc_hd__clkbuf_1 _442_ (.A(_099_),
    .X(_108_));
 sky130_fd_sc_hd__clkbuf_1 _443_ (.A(\mem_top_track_0.DFF_2_.Q ),
    .X(_100_));
 sky130_fd_sc_hd__clkbuf_1 _444_ (.A(_100_),
    .X(_106_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .Y(_118_));
 sky130_fd_sc_hd__clkbuf_1 _446_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_1 _447_ (.A(_101_),
    .X(_109_));
 sky130_fd_sc_hd__clkbuf_1 _448_ (.A(\mem_top_track_0.DFF_2_.Q ),
    .X(_102_));
 sky130_fd_sc_hd__clkbuf_1 _449_ (.A(_102_),
    .X(_105_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .Y(_116_));
 sky130_fd_sc_hd__clkbuf_1 _451_ (.A(\mem_top_track_0.DFF_1_.Q ),
    .X(_103_));
 sky130_fd_sc_hd__clkbuf_1 _452_ (.A(_103_),
    .X(_107_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(\mux_top_track_0.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _454_ (.A(net44),
    .Y(\mux_top_track_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _455_ (.A(\mux_top_track_8.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _456_ (.A(net45),
    .Y(\mux_top_track_8.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _457_ (.A(\mux_right_track_0.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _458_ (.A(net43),
    .Y(\mux_right_track_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _459_ (.A(\mux_right_track_8.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _460_ (.A(net42),
    .Y(\mux_right_track_8.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _461_ (.A(\mux_bottom_track_1.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net65));
 sky130_fd_sc_hd__inv_2 _462_ (.A(net9),
    .Y(\mux_bottom_track_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _463_ (.A(net5),
    .Y(\mux_bottom_track_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _464_ (.A(net2),
    .Y(\mux_bottom_track_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _465_ (.A(net20),
    .Y(\mux_bottom_track_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _466_ (.A(net18),
    .Y(\mux_bottom_track_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _467_ (.A(net14),
    .Y(\mux_bottom_track_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _468_ (.A(net35),
    .Y(\mux_bottom_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _469_ (.A(net31),
    .Y(\mux_bottom_track_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _470_ (.A(net11),
    .Y(\mux_bottom_track_1.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _471_ (.A(\mux_bottom_track_9.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _472_ (.A(net10),
    .Y(\mux_bottom_track_9.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _473_ (.A(net6),
    .Y(\mux_bottom_track_9.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _474_ (.A(net1),
    .Y(\mux_bottom_track_9.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _475_ (.A(net17),
    .Y(\mux_bottom_track_9.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _476_ (.A(net16),
    .Y(\mux_bottom_track_9.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _477_ (.A(net13),
    .Y(\mux_bottom_track_9.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _478_ (.A(net36),
    .Y(\mux_bottom_track_9.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _479_ (.A(net32),
    .Y(\mux_bottom_track_9.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _480_ (.A(net12),
    .Y(\mux_bottom_track_9.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _481_ (.A(\mux_left_track_1.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net47));
 sky130_fd_sc_hd__inv_2 _482_ (.A(net30),
    .Y(\mux_left_track_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _483_ (.A(net28),
    .Y(\mux_left_track_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _484_ (.A(net24),
    .Y(\mux_left_track_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _485_ (.A(net34),
    .Y(\mux_left_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _486_ (.A(net41),
    .Y(\mux_left_track_1.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _487_ (.A(\mux_left_track_9.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net51));
 sky130_fd_sc_hd__inv_2 _488_ (.A(net26),
    .Y(\mux_left_track_9.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _489_ (.A(net25),
    .Y(\mux_left_track_9.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _490_ (.A(net22),
    .Y(\mux_left_track_9.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _491_ (.A(net39),
    .Y(\mux_left_track_9.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _492_ (.A(net40),
    .Y(\mux_left_track_9.INVTX1_8_.out ));
 sky130_fd_sc_hd__inv_2 _493_ (.A(\mux_top_track_16.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _494_ (.A(\mux_right_track_16.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _495_ (.A(\mux_bottom_track_17.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _496_ (.A(net7),
    .Y(\mux_bottom_track_17.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _497_ (.A(net4),
    .Y(\mux_bottom_track_17.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _498_ (.A(net21),
    .Y(\mux_bottom_track_17.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _499_ (.A(net19),
    .Y(\mux_bottom_track_17.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _500_ (.A(net15),
    .Y(\mux_bottom_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _501_ (.A(net37),
    .Y(\mux_bottom_track_17.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _502_ (.A(net33),
    .Y(\mux_bottom_track_17.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _503_ (.A(net8),
    .Y(\mux_bottom_track_17.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _504_ (.A(\mux_left_track_17.mux_l4_in_0_.TGATE_0_.out ),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _505_ (.A(net27),
    .Y(\mux_left_track_17.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _506_ (.A(net23),
    .Y(\mux_left_track_17.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _507_ (.A(net38),
    .Y(\mux_left_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _508_ (.A(net29),
    .Y(\mux_left_track_17.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _509_ (.A(net46),
    .Y(_304_));
 sky130_fd_sc_hd__inv_2 _510_ (.A(\mem_left_track_17.DFF_2_.Q ),
    .Y(_306_));
 sky130_fd_sc_hd__inv_2 _511_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .Y(_310_));
 sky130_fd_sc_hd__inv_2 _512_ (.A(\mem_left_track_17.DFF_0_.Q ),
    .Y(_311_));
 sky130_fd_sc_hd__clkbuf_1 _513_ (.A(\mem_top_track_0.DFF_3_.Q ),
    .X(_000_));
 sky130_fd_sc_hd__clkbuf_1 _514_ (.A(_000_),
    .X(_104_));
 sky130_fd_sc_hd__clkbuf_1 _515_ (.A(\mem_left_track_17.DFF_0_.Q ),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_1 _516_ (.A(_001_),
    .X(_303_));
 sky130_fd_sc_hd__clkbuf_1 _517_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .X(_002_));
 sky130_fd_sc_hd__clkbuf_1 _518_ (.A(_002_),
    .X(_302_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(\mem_left_track_17.DFF_2_.Q ),
    .X(_003_));
 sky130_fd_sc_hd__clkbuf_1 _520_ (.A(_003_),
    .X(_298_));
 sky130_fd_sc_hd__inv_2 _521_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .Y(_309_));
 sky130_fd_sc_hd__clkbuf_1 _522_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .X(_004_));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(_004_),
    .X(_301_));
 sky130_fd_sc_hd__clkbuf_1 _524_ (.A(net46),
    .X(_005_));
 sky130_fd_sc_hd__buf_1 _525_ (.A(_005_),
    .X(_296_));
 sky130_fd_sc_hd__inv_2 _526_ (.A(\mem_left_track_17.DFF_2_.Q ),
    .Y(_305_));
 sky130_fd_sc_hd__inv_2 _527_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .Y(_308_));
 sky130_fd_sc_hd__clkbuf_1 _528_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .X(_006_));
 sky130_fd_sc_hd__clkbuf_1 _529_ (.A(_006_),
    .X(_300_));
 sky130_fd_sc_hd__clkbuf_1 _530_ (.A(\mem_left_track_17.DFF_2_.Q ),
    .X(_007_));
 sky130_fd_sc_hd__clkbuf_1 _531_ (.A(_007_),
    .X(_297_));
 sky130_fd_sc_hd__inv_2 _532_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .Y(_307_));
 sky130_fd_sc_hd__clkbuf_1 _533_ (.A(\mem_left_track_17.DFF_1_.Q ),
    .X(_008_));
 sky130_fd_sc_hd__clkbuf_1 _534_ (.A(_008_),
    .X(_299_));
 sky130_fd_sc_hd__inv_2 _535_ (.A(\mem_bottom_track_17.DFF_3_.Q ),
    .Y(_288_));
 sky130_fd_sc_hd__inv_2 _536_ (.A(\mem_bottom_track_17.DFF_2_.Q ),
    .Y(_290_));
 sky130_fd_sc_hd__inv_2 _537_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .Y(_294_));
 sky130_fd_sc_hd__inv_2 _538_ (.A(\mem_bottom_track_17.DFF_0_.Q ),
    .Y(_295_));
 sky130_fd_sc_hd__clkbuf_1 _539_ (.A(\mem_bottom_track_17.DFF_0_.Q ),
    .X(_009_));
 sky130_fd_sc_hd__clkbuf_1 _540_ (.A(_009_),
    .X(_287_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .X(_010_));
 sky130_fd_sc_hd__clkbuf_1 _542_ (.A(_010_),
    .X(_286_));
 sky130_fd_sc_hd__clkbuf_1 _543_ (.A(\mem_bottom_track_17.DFF_2_.Q ),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_1 _544_ (.A(_011_),
    .X(_282_));
 sky130_fd_sc_hd__inv_2 _545_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .Y(_293_));
 sky130_fd_sc_hd__clkbuf_1 _546_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .X(_012_));
 sky130_fd_sc_hd__clkbuf_1 _547_ (.A(_012_),
    .X(_285_));
 sky130_fd_sc_hd__clkbuf_1 _548_ (.A(\mem_bottom_track_17.DFF_3_.Q ),
    .X(_013_));
 sky130_fd_sc_hd__clkbuf_1 _549_ (.A(_013_),
    .X(_280_));
 sky130_fd_sc_hd__inv_2 _550_ (.A(\mem_bottom_track_17.DFF_2_.Q ),
    .Y(_289_));
 sky130_fd_sc_hd__inv_2 _551_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .Y(_292_));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .X(_014_));
 sky130_fd_sc_hd__clkbuf_1 _553_ (.A(_014_),
    .X(_284_));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(\mem_bottom_track_17.DFF_2_.Q ),
    .X(_015_));
 sky130_fd_sc_hd__clkbuf_1 _555_ (.A(_015_),
    .X(_281_));
 sky130_fd_sc_hd__inv_2 _556_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .Y(_291_));
 sky130_fd_sc_hd__clkbuf_1 _557_ (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .X(_016_));
 sky130_fd_sc_hd__clkbuf_1 _558_ (.A(_016_),
    .X(_283_));
 sky130_fd_sc_hd__inv_2 _559_ (.A(\mem_bottom_track_1.DFF_0_.D ),
    .Y(_272_));
 sky130_fd_sc_hd__inv_2 _560_ (.A(\mem_right_track_16.DFF_2_.Q ),
    .Y(_274_));
 sky130_fd_sc_hd__inv_2 _561_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .Y(_278_));
 sky130_fd_sc_hd__inv_2 _562_ (.A(\mem_right_track_16.DFF_0_.Q ),
    .Y(_279_));
 sky130_fd_sc_hd__clkbuf_1 _563_ (.A(\mem_right_track_16.DFF_0_.Q ),
    .X(_017_));
 sky130_fd_sc_hd__clkbuf_1 _564_ (.A(_017_),
    .X(_271_));
 sky130_fd_sc_hd__clkbuf_1 _565_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .X(_018_));
 sky130_fd_sc_hd__clkbuf_1 _566_ (.A(_018_),
    .X(_270_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(\mem_right_track_16.DFF_2_.Q ),
    .X(_019_));
 sky130_fd_sc_hd__clkbuf_1 _568_ (.A(_019_),
    .X(_266_));
 sky130_fd_sc_hd__inv_2 _569_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .Y(_277_));
 sky130_fd_sc_hd__clkbuf_1 _570_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .X(_020_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_020_),
    .X(_269_));
 sky130_fd_sc_hd__clkbuf_1 _572_ (.A(\mem_bottom_track_1.DFF_0_.D ),
    .X(_021_));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(_021_),
    .X(_264_));
 sky130_fd_sc_hd__inv_2 _574_ (.A(\mem_right_track_16.DFF_2_.Q ),
    .Y(_273_));
 sky130_fd_sc_hd__inv_2 _575_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .Y(_276_));
 sky130_fd_sc_hd__clkbuf_1 _576_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .X(_022_));
 sky130_fd_sc_hd__clkbuf_1 _577_ (.A(_022_),
    .X(_268_));
 sky130_fd_sc_hd__clkbuf_1 _578_ (.A(\mem_right_track_16.DFF_2_.Q ),
    .X(_023_));
 sky130_fd_sc_hd__clkbuf_1 _579_ (.A(_023_),
    .X(_265_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .Y(_275_));
 sky130_fd_sc_hd__clkbuf_1 _581_ (.A(\mem_right_track_16.DFF_1_.Q ),
    .X(_024_));
 sky130_fd_sc_hd__clkbuf_1 _582_ (.A(_024_),
    .X(_267_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(\mem_right_track_0.DFF_0_.D ),
    .Y(_256_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(\mem_top_track_16.DFF_2_.Q ),
    .Y(_258_));
 sky130_fd_sc_hd__inv_2 _585_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .Y(_262_));
 sky130_fd_sc_hd__inv_2 _586_ (.A(\mem_top_track_16.DFF_0_.Q ),
    .Y(_263_));
 sky130_fd_sc_hd__clkbuf_1 _587_ (.A(\mem_top_track_16.DFF_0_.Q ),
    .X(_025_));
 sky130_fd_sc_hd__clkbuf_1 _588_ (.A(_025_),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _589_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .X(_026_));
 sky130_fd_sc_hd__clkbuf_1 _590_ (.A(_026_),
    .X(_254_));
 sky130_fd_sc_hd__clkbuf_1 _591_ (.A(\mem_top_track_16.DFF_2_.Q ),
    .X(_027_));
 sky130_fd_sc_hd__clkbuf_1 _592_ (.A(_027_),
    .X(_250_));
 sky130_fd_sc_hd__inv_2 _593_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .Y(_261_));
 sky130_fd_sc_hd__clkbuf_1 _594_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .X(_028_));
 sky130_fd_sc_hd__clkbuf_1 _595_ (.A(_028_),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _596_ (.A(\mem_right_track_0.DFF_0_.D ),
    .X(_029_));
 sky130_fd_sc_hd__clkbuf_1 _597_ (.A(_029_),
    .X(_248_));
 sky130_fd_sc_hd__inv_2 _598_ (.A(\mem_top_track_16.DFF_2_.Q ),
    .Y(_257_));
 sky130_fd_sc_hd__inv_2 _599_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .Y(_260_));
 sky130_fd_sc_hd__clkbuf_1 _600_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .X(_030_));
 sky130_fd_sc_hd__clkbuf_1 _601_ (.A(_030_),
    .X(_252_));
 sky130_fd_sc_hd__clkbuf_1 _602_ (.A(\mem_top_track_16.DFF_2_.Q ),
    .X(_031_));
 sky130_fd_sc_hd__clkbuf_1 _603_ (.A(_031_),
    .X(_249_));
 sky130_fd_sc_hd__inv_2 _604_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .Y(_259_));
 sky130_fd_sc_hd__clkbuf_1 _605_ (.A(\mem_top_track_16.DFF_1_.Q ),
    .X(_032_));
 sky130_fd_sc_hd__clkbuf_1 _606_ (.A(_032_),
    .X(_251_));
 sky130_fd_sc_hd__inv_2 _607_ (.A(\mem_left_track_17.DFF_0_.D ),
    .Y(_239_));
 sky130_fd_sc_hd__inv_2 _608_ (.A(\mem_left_track_9.DFF_2_.Q ),
    .Y(_241_));
 sky130_fd_sc_hd__inv_2 _609_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .Y(_245_));
 sky130_fd_sc_hd__inv_2 _610_ (.A(\mem_left_track_9.DFF_0_.Q ),
    .Y(_247_));
 sky130_fd_sc_hd__clkbuf_1 _611_ (.A(\mem_left_track_9.DFF_0_.Q ),
    .X(_033_));
 sky130_fd_sc_hd__clkbuf_1 _612_ (.A(_033_),
    .X(_238_));
 sky130_fd_sc_hd__clkbuf_1 _613_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_1 _614_ (.A(_034_),
    .X(_236_));
 sky130_fd_sc_hd__inv_2 _615_ (.A(\mem_left_track_9.DFF_0_.Q ),
    .Y(_246_));
 sky130_fd_sc_hd__clkbuf_1 _616_ (.A(\mem_left_track_9.DFF_0_.Q ),
    .X(_035_));
 sky130_fd_sc_hd__clkbuf_1 _617_ (.A(_035_),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _618_ (.A(\mem_left_track_9.DFF_2_.Q ),
    .X(_036_));
 sky130_fd_sc_hd__clkbuf_1 _619_ (.A(_036_),
    .X(_232_));
 sky130_fd_sc_hd__inv_2 _620_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .Y(_244_));
 sky130_fd_sc_hd__clkbuf_1 _621_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .X(_037_));
 sky130_fd_sc_hd__clkbuf_1 _622_ (.A(_037_),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _623_ (.A(\mem_left_track_17.DFF_0_.D ),
    .X(_038_));
 sky130_fd_sc_hd__clkbuf_1 _624_ (.A(_038_),
    .X(_230_));
 sky130_fd_sc_hd__inv_2 _625_ (.A(\mem_left_track_9.DFF_2_.Q ),
    .Y(_240_));
 sky130_fd_sc_hd__inv_2 _626_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .Y(_243_));
 sky130_fd_sc_hd__clkbuf_1 _627_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .X(_039_));
 sky130_fd_sc_hd__clkbuf_1 _628_ (.A(_039_),
    .X(_234_));
 sky130_fd_sc_hd__clkbuf_1 _629_ (.A(\mem_left_track_9.DFF_2_.Q ),
    .X(_040_));
 sky130_fd_sc_hd__clkbuf_1 _630_ (.A(_040_),
    .X(_231_));
 sky130_fd_sc_hd__inv_2 _631_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .Y(_242_));
 sky130_fd_sc_hd__clkbuf_1 _632_ (.A(\mem_left_track_9.DFF_1_.Q ),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_1 _633_ (.A(_041_),
    .X(_233_));
 sky130_fd_sc_hd__inv_2 _634_ (.A(\mem_left_track_1.DFF_3_.Q ),
    .Y(_221_));
 sky130_fd_sc_hd__inv_2 _635_ (.A(\mem_left_track_1.DFF_2_.Q ),
    .Y(_223_));
 sky130_fd_sc_hd__inv_2 _636_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .Y(_227_));
 sky130_fd_sc_hd__inv_2 _637_ (.A(\mem_left_track_1.DFF_0_.Q ),
    .Y(_229_));
 sky130_fd_sc_hd__clkbuf_1 _638_ (.A(\mem_left_track_1.DFF_0_.Q ),
    .X(_042_));
 sky130_fd_sc_hd__clkbuf_1 _639_ (.A(_042_),
    .X(_220_));
 sky130_fd_sc_hd__clkbuf_1 _640_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .X(_043_));
 sky130_fd_sc_hd__clkbuf_1 _641_ (.A(_043_),
    .X(_218_));
 sky130_fd_sc_hd__inv_2 _642_ (.A(\mem_left_track_1.DFF_0_.Q ),
    .Y(_228_));
 sky130_fd_sc_hd__clkbuf_1 _643_ (.A(\mem_left_track_1.DFF_0_.Q ),
    .X(_044_));
 sky130_fd_sc_hd__clkbuf_1 _644_ (.A(_044_),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_1 _645_ (.A(\mem_left_track_1.DFF_2_.Q ),
    .X(_045_));
 sky130_fd_sc_hd__clkbuf_1 _646_ (.A(_045_),
    .X(_214_));
 sky130_fd_sc_hd__inv_2 _647_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .Y(_226_));
 sky130_fd_sc_hd__clkbuf_1 _648_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .X(_046_));
 sky130_fd_sc_hd__clkbuf_1 _649_ (.A(_046_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _650_ (.A(\mem_left_track_1.DFF_3_.Q ),
    .X(_047_));
 sky130_fd_sc_hd__clkbuf_1 _651_ (.A(_047_),
    .X(_212_));
 sky130_fd_sc_hd__inv_2 _652_ (.A(\mem_left_track_1.DFF_2_.Q ),
    .Y(_222_));
 sky130_fd_sc_hd__inv_2 _653_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .Y(_225_));
 sky130_fd_sc_hd__clkbuf_1 _654_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _655_ (.A(_048_),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _656_ (.A(\mem_left_track_1.DFF_2_.Q ),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _657_ (.A(_049_),
    .X(_213_));
 sky130_fd_sc_hd__inv_2 _658_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .Y(_224_));
 sky130_fd_sc_hd__clkbuf_1 _659_ (.A(\mem_left_track_1.DFF_1_.Q ),
    .X(_050_));
 sky130_fd_sc_hd__clkbuf_1 _660_ (.A(_050_),
    .X(_215_));
 sky130_fd_sc_hd__inv_2 _661_ (.A(\mem_bottom_track_17.DFF_0_.D ),
    .Y(_203_));
 sky130_fd_sc_hd__inv_2 _662_ (.A(\mem_bottom_track_9.DFF_2_.Q ),
    .Y(_205_));
 sky130_fd_sc_hd__inv_2 _663_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .Y(_209_));
 sky130_fd_sc_hd__inv_2 _664_ (.A(\mem_bottom_track_9.DFF_0_.Q ),
    .Y(_211_));
 sky130_fd_sc_hd__clkbuf_1 _665_ (.A(\mem_bottom_track_9.DFF_0_.Q ),
    .X(_051_));
 sky130_fd_sc_hd__clkbuf_1 _666_ (.A(_051_),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _667_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .X(_052_));
 sky130_fd_sc_hd__clkbuf_1 _668_ (.A(_052_),
    .X(_200_));
 sky130_fd_sc_hd__inv_2 _669_ (.A(\mem_bottom_track_9.DFF_0_.Q ),
    .Y(_210_));
 sky130_fd_sc_hd__clkbuf_1 _670_ (.A(\mem_bottom_track_9.DFF_0_.Q ),
    .X(_053_));
 sky130_fd_sc_hd__clkbuf_1 _671_ (.A(_053_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _672_ (.A(\mem_bottom_track_9.DFF_2_.Q ),
    .X(_054_));
 sky130_fd_sc_hd__clkbuf_1 _673_ (.A(_054_),
    .X(_196_));
 sky130_fd_sc_hd__inv_2 _674_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .Y(_208_));
 sky130_fd_sc_hd__clkbuf_1 _675_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .X(_055_));
 sky130_fd_sc_hd__clkbuf_1 _676_ (.A(_055_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _677_ (.A(\mem_bottom_track_17.DFF_0_.D ),
    .X(_056_));
 sky130_fd_sc_hd__clkbuf_1 _678_ (.A(_056_),
    .X(_194_));
 sky130_fd_sc_hd__inv_2 _679_ (.A(\mem_bottom_track_9.DFF_2_.Q ),
    .Y(_204_));
 sky130_fd_sc_hd__inv_2 _680_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .Y(_207_));
 sky130_fd_sc_hd__clkbuf_1 _681_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .X(_057_));
 sky130_fd_sc_hd__clkbuf_1 _682_ (.A(_057_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _683_ (.A(\mem_bottom_track_9.DFF_2_.Q ),
    .X(_058_));
 sky130_fd_sc_hd__clkbuf_1 _684_ (.A(_058_),
    .X(_195_));
 sky130_fd_sc_hd__inv_2 _685_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .Y(_206_));
 sky130_fd_sc_hd__clkbuf_1 _686_ (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .X(_059_));
 sky130_fd_sc_hd__clkbuf_1 _687_ (.A(_059_),
    .X(_197_));
 sky130_fd_sc_hd__inv_2 _688_ (.A(\mem_bottom_track_1.DFF_3_.Q ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_2 _689_ (.A(\mem_bottom_track_1.DFF_2_.Q ),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _690_ (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .Y(_191_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(\mem_bottom_track_1.DFF_0_.Q ),
    .Y(_193_));
 sky130_fd_sc_hd__dfxtp_1 _692_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net118),
    .Q(\mem_top_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _693_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net139),
    .Q(\mem_top_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _694_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net126),
    .Q(\mem_top_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _695_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net3),
    .Q(\mem_top_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _696_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net127),
    .Q(\mem_top_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _697_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net135),
    .Q(\mem_top_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _698_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net110),
    .Q(\mem_top_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _699_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net106),
    .Q(\mem_top_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _700_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net117),
    .Q(\mem_right_track_0.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _701_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net131),
    .Q(\mem_right_track_0.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _702_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net128),
    .Q(\mem_right_track_0.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _703_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net96),
    .Q(\mem_right_track_0.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _704_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net116),
    .Q(\mem_right_track_16.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _705_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net132),
    .Q(\mem_right_track_8.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _706_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net113),
    .Q(\mem_right_track_8.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _707_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net103),
    .Q(\mem_right_track_8.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _708_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net119),
    .Q(\mem_bottom_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _709_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net137),
    .Q(\mem_bottom_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _710_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net111),
    .Q(\mem_bottom_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _711_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net95),
    .Q(\mem_bottom_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _712_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net115),
    .Q(\mem_bottom_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _713_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net123),
    .Q(\mem_bottom_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _714_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net130),
    .Q(\mem_bottom_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _715_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net98),
    .Q(\mem_bottom_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _716_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net121),
    .Q(\mem_left_track_1.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _717_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net133),
    .Q(\mem_left_track_1.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _718_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net109),
    .Q(\mem_left_track_1.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _719_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net105),
    .Q(\mem_left_track_1.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _720_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net122),
    .Q(\mem_left_track_17.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _721_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net140),
    .Q(\mem_left_track_9.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _722_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net120),
    .Q(\mem_left_track_9.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _723_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net108),
    .Q(\mem_left_track_9.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _724_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net125),
    .Q(\mem_right_track_0.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _725_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net138),
    .Q(\mem_top_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _726_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net97),
    .Q(\mem_top_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _727_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net104),
    .Q(\mem_top_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _728_ (.CLK(clknet_2_0__leaf_prog_clk),
    .D(net114),
    .Q(\mem_bottom_track_1.DFF_0_.D ));
 sky130_fd_sc_hd__dfxtp_1 _729_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net141),
    .Q(\mem_right_track_16.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _730_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net100),
    .Q(\mem_right_track_16.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _731_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net101),
    .Q(\mem_right_track_16.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _732_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net129),
    .Q(\mem_bottom_track_17.DFF_3_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _733_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net134),
    .Q(\mem_bottom_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _734_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net112),
    .Q(\mem_bottom_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _735_ (.CLK(clknet_2_1__leaf_prog_clk),
    .D(net102),
    .Q(\mem_bottom_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _736_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net124),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_2 _737_ (.CLK(clknet_2_3__leaf_prog_clk),
    .D(net136),
    .Q(\mem_left_track_17.DFF_2_.Q ));
 sky130_fd_sc_hd__dfxtp_2 _738_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net107),
    .Q(\mem_left_track_17.DFF_1_.Q ));
 sky130_fd_sc_hd__dfxtp_1 _739_ (.CLK(clknet_2_2__leaf_prog_clk),
    .D(net99),
    .Q(\mem_left_track_17.DFF_0_.Q ));
 sky130_fd_sc_hd__buf_1 _752_ (.A(net19),
    .X(net54));
 sky130_fd_sc_hd__buf_1 _753_ (.A(net18),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _754_ (.A(net17),
    .X(net52));
 sky130_fd_sc_hd__buf_1 _755_ (.A(net15),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _756_ (.A(net14),
    .X(net49));
 sky130_fd_sc_hd__buf_1 _757_ (.A(net13),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _758_ (.A(net10),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _759_ (.A(net9),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _760_ (.A(net8),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _761_ (.A(net6),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _762_ (.A(net5),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _763_ (.A(net4),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _764_ (.A(net37),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 _765_ (.A(net36),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _766_ (.A(net35),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _767_ (.A(net33),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _768_ (.A(net32),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _769_ (.A(net31),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _770_ (.A(net28),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _771_ (.A(net27),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _772_ (.A(net26),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _773_ (.A(net24),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _774_ (.A(net23),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _775_ (.A(net22),
    .X(net75));
 sky130_fd_sc_hd__ebufn_2 _776_ (.A(\mux_top_track_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_104_),
    .Z(\mux_top_track_0.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _777_ (.A(\mux_top_track_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_105_),
    .Z(\mux_top_track_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _778_ (.A(\mux_top_track_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_106_),
    .Z(\mux_top_track_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _779_ (.A(net83),
    .TE_B(_107_),
    .Z(\mux_top_track_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _779__83 (.HI(net83));
 sky130_fd_sc_hd__ebufn_1 _780_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_108_),
    .Z(\mux_top_track_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _781_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_109_),
    .Z(\mux_top_track_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _782_ (.A(\mux_top_track_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_110_),
    .Z(\mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _783_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_111_),
    .Z(\mux_top_track_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _784_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_112_),
    .Z(\mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _785_ (.A(\mux_top_track_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_113_),
    .Z(\mux_top_track_0.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _786_ (.A(\mux_top_track_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_114_),
    .Z(\mux_top_track_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _787_ (.A(\mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_115_),
    .Z(\mux_top_track_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _788_ (.A(\mux_bottom_track_17.INVTX1_7_.out ),
    .TE_B(_116_),
    .Z(\mux_top_track_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _789_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_117_),
    .Z(\mux_top_track_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _790_ (.A(\mux_left_track_9.INVTX1_5_.out ),
    .TE_B(_118_),
    .Z(\mux_top_track_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _791_ (.A(\mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_119_),
    .Z(\mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _792_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_120_),
    .Z(\mux_top_track_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _793_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_121_),
    .Z(\mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _794_ (.A(\mux_top_track_8.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_122_),
    .Z(\mux_top_track_8.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _795_ (.A(\mux_top_track_8.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_123_),
    .Z(\mux_top_track_8.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _796_ (.A(\mux_top_track_8.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_124_),
    .Z(\mux_top_track_8.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _797_ (.A(net84),
    .TE_B(_125_),
    .Z(\mux_top_track_8.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _797__84 (.HI(net84));
 sky130_fd_sc_hd__ebufn_1 _798_ (.A(\mux_bottom_track_9.INVTX1_7_.out ),
    .TE_B(_126_),
    .Z(\mux_top_track_8.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _799_ (.A(\mux_left_track_17.INVTX1_6_.out ),
    .TE_B(_127_),
    .Z(\mux_top_track_8.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _800_ (.A(\mux_top_track_8.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_128_),
    .Z(\mux_top_track_8.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _801_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_129_),
    .Z(\mux_top_track_8.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _802_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_130_),
    .Z(\mux_top_track_8.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _803_ (.A(\mux_top_track_8.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_131_),
    .Z(\mux_top_track_8.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _804_ (.A(\mux_top_track_8.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_132_),
    .Z(\mux_top_track_8.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _805_ (.A(\mux_top_track_8.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_133_),
    .Z(\mux_top_track_8.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _806_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_134_),
    .Z(\mux_top_track_8.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _807_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_135_),
    .Z(\mux_top_track_8.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _808_ (.A(\mux_left_track_17.INVTX1_5_.out ),
    .TE_B(_136_),
    .Z(\mux_top_track_8.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _809_ (.A(\mux_top_track_8.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_137_),
    .Z(\mux_top_track_8.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _810_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_138_),
    .Z(\mux_top_track_8.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _811_ (.A(\mux_top_track_8.INVTX1_0_.out ),
    .TE_B(_139_),
    .Z(\mux_top_track_8.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _812_ (.A(\mux_right_track_0.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_140_),
    .Z(\mux_right_track_0.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _813_ (.A(\mux_right_track_0.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_141_),
    .Z(\mux_right_track_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _814_ (.A(\mux_right_track_0.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_142_),
    .Z(\mux_right_track_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _815_ (.A(net85),
    .TE_B(_143_),
    .Z(\mux_right_track_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _815__85 (.HI(net85));
 sky130_fd_sc_hd__ebufn_1 _816_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_144_),
    .Z(\mux_right_track_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _817_ (.A(\mux_left_track_17.INVTX1_6_.out ),
    .TE_B(_145_),
    .Z(\mux_right_track_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _818_ (.A(\mux_right_track_0.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_146_),
    .Z(\mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _819_ (.A(\mux_right_track_0.INVTX1_3_.out ),
    .TE_B(_147_),
    .Z(\mux_right_track_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _820_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_148_),
    .Z(\mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _821_ (.A(\mux_right_track_0.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_149_),
    .Z(\mux_right_track_0.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _822_ (.A(\mux_right_track_0.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_150_),
    .Z(\mux_right_track_0.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _823_ (.A(\mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_151_),
    .Z(\mux_right_track_0.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _824_ (.A(\mux_bottom_track_17.INVTX1_7_.out ),
    .TE_B(_152_),
    .Z(\mux_right_track_0.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _825_ (.A(\mux_left_track_17.INVTX1_7_.out ),
    .TE_B(_153_),
    .Z(\mux_right_track_0.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _826_ (.A(\mux_left_track_17.INVTX1_5_.out ),
    .TE_B(_154_),
    .Z(\mux_right_track_0.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _827_ (.A(\mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_155_),
    .Z(\mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _828_ (.A(\mux_left_track_9.INVTX1_2_.out ),
    .TE_B(_156_),
    .Z(\mux_right_track_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _829_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_157_),
    .Z(\mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _830_ (.A(\mux_right_track_8.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_158_),
    .Z(\mux_right_track_8.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _831_ (.A(\mux_right_track_8.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_159_),
    .Z(\mux_right_track_8.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _832_ (.A(\mux_right_track_8.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_160_),
    .Z(\mux_right_track_8.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _833_ (.A(net86),
    .TE_B(_161_),
    .Z(\mux_right_track_8.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _833__86 (.HI(net86));
 sky130_fd_sc_hd__ebufn_1 _834_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_162_),
    .Z(\mux_right_track_8.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _835_ (.A(\mux_left_track_9.INVTX1_6_.out ),
    .TE_B(_163_),
    .Z(\mux_right_track_8.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _836_ (.A(\mux_right_track_8.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_164_),
    .Z(\mux_right_track_8.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _837_ (.A(\mux_right_track_8.INVTX1_3_.out ),
    .TE_B(_165_),
    .Z(\mux_right_track_8.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _838_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_166_),
    .Z(\mux_right_track_8.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _839_ (.A(\mux_right_track_8.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_167_),
    .Z(\mux_right_track_8.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _840_ (.A(\mux_right_track_8.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_168_),
    .Z(\mux_right_track_8.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _841_ (.A(\mux_right_track_8.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_169_),
    .Z(\mux_right_track_8.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _842_ (.A(\mux_bottom_track_1.INVTX1_7_.out ),
    .TE_B(_170_),
    .Z(\mux_right_track_8.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _843_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_171_),
    .Z(\mux_right_track_8.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _844_ (.A(\mux_left_track_9.INVTX1_5_.out ),
    .TE_B(_172_),
    .Z(\mux_right_track_8.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _845_ (.A(\mux_right_track_8.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_173_),
    .Z(\mux_right_track_8.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _846_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_174_),
    .Z(\mux_right_track_8.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _847_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_175_),
    .Z(\mux_right_track_8.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _848_ (.A(\mux_bottom_track_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_176_),
    .Z(\mux_bottom_track_1.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _849_ (.A(\mux_bottom_track_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_177_),
    .Z(\mux_bottom_track_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _850_ (.A(\mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_178_),
    .Z(\mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _851_ (.A(net87),
    .TE_B(_179_),
    .Z(\mux_bottom_track_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _851__87 (.HI(net87));
 sky130_fd_sc_hd__ebufn_1 _852_ (.A(\mux_bottom_track_1.INVTX1_7_.out ),
    .TE_B(_180_),
    .Z(\mux_bottom_track_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _853_ (.A(\mux_bottom_track_1.INVTX1_5_.out ),
    .TE_B(_181_),
    .Z(\mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _854_ (.A(\mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_182_),
    .Z(\mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _855_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_183_),
    .Z(\mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _856_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_184_),
    .Z(\mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _857_ (.A(\mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_185_),
    .Z(\mux_bottom_track_1.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _858_ (.A(\mux_bottom_track_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_186_),
    .Z(\mux_bottom_track_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _859_ (.A(\mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_187_),
    .Z(\mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _860_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_188_),
    .Z(\mux_bottom_track_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _861_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_189_),
    .Z(\mux_bottom_track_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _862_ (.A(\mux_bottom_track_1.INVTX1_4_.out ),
    .TE_B(_190_),
    .Z(\mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _863_ (.A(\mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_191_),
    .Z(\mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _864_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_192_),
    .Z(\mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _865_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_193_),
    .Z(\mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _866_ (.A(\mux_bottom_track_9.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_194_),
    .Z(\mux_bottom_track_9.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _867_ (.A(\mux_bottom_track_9.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_195_),
    .Z(\mux_bottom_track_9.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _868_ (.A(\mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_196_),
    .Z(\mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _869_ (.A(net88),
    .TE_B(_197_),
    .Z(\mux_bottom_track_9.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _869__88 (.HI(net88));
 sky130_fd_sc_hd__ebufn_1 _870_ (.A(\mux_bottom_track_9.INVTX1_7_.out ),
    .TE_B(_198_),
    .Z(\mux_bottom_track_9.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _871_ (.A(\mux_bottom_track_9.INVTX1_5_.out ),
    .TE_B(_199_),
    .Z(\mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _872_ (.A(\mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_200_),
    .Z(\mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _873_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_201_),
    .Z(\mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _874_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_202_),
    .Z(\mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _875_ (.A(\mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_203_),
    .Z(\mux_bottom_track_9.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _876_ (.A(\mux_bottom_track_9.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_204_),
    .Z(\mux_bottom_track_9.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _877_ (.A(\mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_205_),
    .Z(\mux_bottom_track_9.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _878_ (.A(\mux_bottom_track_9.INVTX1_8_.out ),
    .TE_B(_206_),
    .Z(\mux_bottom_track_9.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _879_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_207_),
    .Z(\mux_bottom_track_9.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _880_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_208_),
    .Z(\mux_bottom_track_9.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _881_ (.A(\mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_209_),
    .Z(\mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _882_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_210_),
    .Z(\mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _883_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_211_),
    .Z(\mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _884_ (.A(\mux_left_track_1.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_212_),
    .Z(\mux_left_track_1.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _885_ (.A(\mux_left_track_1.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_213_),
    .Z(\mux_left_track_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _886_ (.A(\mux_left_track_1.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_214_),
    .Z(\mux_left_track_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _887_ (.A(net89),
    .TE_B(_215_),
    .Z(\mux_left_track_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _887__89 (.HI(net89));
 sky130_fd_sc_hd__ebufn_1 _888_ (.A(\mux_left_track_1.INVTX1_7_.out ),
    .TE_B(_216_),
    .Z(\mux_left_track_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _889_ (.A(\mux_left_track_1.INVTX1_5_.out ),
    .TE_B(_217_),
    .Z(\mux_left_track_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _890_ (.A(\mux_left_track_1.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_218_),
    .Z(\mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _891_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_219_),
    .Z(\mux_left_track_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _892_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_220_),
    .Z(\mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _893_ (.A(\mux_left_track_1.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_221_),
    .Z(\mux_left_track_1.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _894_ (.A(\mux_left_track_1.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_222_),
    .Z(\mux_left_track_1.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _895_ (.A(\mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_223_),
    .Z(\mux_left_track_1.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _896_ (.A(\mux_left_track_1.INVTX1_8_.out ),
    .TE_B(_224_),
    .Z(\mux_left_track_1.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _897_ (.A(\mux_left_track_1.INVTX1_6_.out ),
    .TE_B(_225_),
    .Z(\mux_left_track_1.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _898_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_226_),
    .Z(\mux_left_track_1.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _899_ (.A(\mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_227_),
    .Z(\mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _900_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_228_),
    .Z(\mux_left_track_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _901_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_229_),
    .Z(\mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _902_ (.A(\mux_left_track_9.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_230_),
    .Z(\mux_left_track_9.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _903_ (.A(\mux_left_track_9.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_231_),
    .Z(\mux_left_track_9.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _904_ (.A(\mux_left_track_9.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_232_),
    .Z(\mux_left_track_9.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _905_ (.A(net90),
    .TE_B(_233_),
    .Z(\mux_left_track_9.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _905__90 (.HI(net90));
 sky130_fd_sc_hd__ebufn_1 _906_ (.A(\mux_left_track_9.INVTX1_7_.out ),
    .TE_B(_234_),
    .Z(\mux_left_track_9.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _907_ (.A(\mux_left_track_9.INVTX1_5_.out ),
    .TE_B(_235_),
    .Z(\mux_left_track_9.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _908_ (.A(\mux_left_track_9.mux_l1_in_1_.TGATE_0_.out ),
    .TE_B(_236_),
    .Z(\mux_left_track_9.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _909_ (.A(\mux_bottom_track_1.INVTX1_2_.out ),
    .TE_B(_237_),
    .Z(\mux_left_track_9.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _910_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_238_),
    .Z(\mux_left_track_9.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _911_ (.A(\mux_left_track_9.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_239_),
    .Z(\mux_left_track_9.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _912_ (.A(\mux_left_track_9.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_240_),
    .Z(\mux_left_track_9.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _913_ (.A(\mux_left_track_9.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_241_),
    .Z(\mux_left_track_9.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _914_ (.A(\mux_left_track_9.INVTX1_8_.out ),
    .TE_B(_242_),
    .Z(\mux_left_track_9.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _915_ (.A(\mux_left_track_9.INVTX1_6_.out ),
    .TE_B(_243_),
    .Z(\mux_left_track_9.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _916_ (.A(\mux_bottom_track_1.INVTX1_3_.out ),
    .TE_B(_244_),
    .Z(\mux_left_track_9.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _917_ (.A(\mux_left_track_9.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_245_),
    .Z(\mux_left_track_9.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _918_ (.A(\mux_left_track_9.INVTX1_2_.out ),
    .TE_B(_246_),
    .Z(\mux_left_track_9.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _919_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_247_),
    .Z(\mux_left_track_9.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _920_ (.A(\mux_top_track_16.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_248_),
    .Z(\mux_top_track_16.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _921_ (.A(\mux_top_track_16.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_249_),
    .Z(\mux_top_track_16.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _922_ (.A(\mux_top_track_16.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_250_),
    .Z(\mux_top_track_16.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _923_ (.A(net91),
    .TE_B(_251_),
    .Z(\mux_top_track_16.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _923__91 (.HI(net91));
 sky130_fd_sc_hd__ebufn_1 _924_ (.A(\mux_bottom_track_1.INVTX1_7_.out ),
    .TE_B(_252_),
    .Z(\mux_top_track_16.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _925_ (.A(\mux_left_track_1.INVTX1_6_.out ),
    .TE_B(_253_),
    .Z(\mux_top_track_16.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _926_ (.A(\mux_bottom_track_9.INVTX1_4_.out ),
    .TE_B(_254_),
    .Z(\mux_top_track_16.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _927_ (.A(\mux_bottom_track_9.INVTX1_3_.out ),
    .TE_B(_255_),
    .Z(\mux_top_track_16.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _928_ (.A(\mux_top_track_16.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_256_),
    .Z(\mux_top_track_16.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _929_ (.A(\mux_top_track_16.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_257_),
    .Z(\mux_top_track_16.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _930_ (.A(\mux_top_track_16.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_258_),
    .Z(\mux_top_track_16.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _931_ (.A(\mux_bottom_track_1.INVTX1_8_.out ),
    .TE_B(_259_),
    .Z(\mux_top_track_16.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _932_ (.A(\mux_bottom_track_1.INVTX1_6_.out ),
    .TE_B(_260_),
    .Z(\mux_top_track_16.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _933_ (.A(\mux_left_track_1.INVTX1_5_.out ),
    .TE_B(_261_),
    .Z(\mux_top_track_16.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _934_ (.A(\mux_top_track_16.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_262_),
    .Z(\mux_top_track_16.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _935_ (.A(\mux_bottom_track_9.INVTX1_2_.out ),
    .TE_B(_263_),
    .Z(\mux_top_track_16.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _936_ (.A(\mux_right_track_16.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_264_),
    .Z(\mux_right_track_16.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _937_ (.A(\mux_right_track_16.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_265_),
    .Z(\mux_right_track_16.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _938_ (.A(\mux_right_track_16.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_266_),
    .Z(\mux_right_track_16.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _939_ (.A(net92),
    .TE_B(_267_),
    .Z(\mux_right_track_16.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _939__92 (.HI(net92));
 sky130_fd_sc_hd__ebufn_1 _940_ (.A(\mux_bottom_track_9.INVTX1_6_.out ),
    .TE_B(_268_),
    .Z(\mux_right_track_16.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _941_ (.A(\mux_left_track_1.INVTX1_6_.out ),
    .TE_B(_269_),
    .Z(\mux_right_track_16.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _942_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_270_),
    .Z(\mux_right_track_16.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _943_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_271_),
    .Z(\mux_right_track_16.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _944_ (.A(\mux_right_track_16.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_272_),
    .Z(\mux_right_track_16.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _945_ (.A(\mux_right_track_16.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_273_),
    .Z(\mux_right_track_16.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _946_ (.A(\mux_right_track_16.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_274_),
    .Z(\mux_right_track_16.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _947_ (.A(\mux_bottom_track_9.INVTX1_7_.out ),
    .TE_B(_275_),
    .Z(\mux_right_track_16.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _948_ (.A(\mux_left_track_1.INVTX1_7_.out ),
    .TE_B(_276_),
    .Z(\mux_right_track_16.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _949_ (.A(\mux_left_track_1.INVTX1_5_.out ),
    .TE_B(_277_),
    .Z(\mux_right_track_16.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _950_ (.A(\mux_right_track_16.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_278_),
    .Z(\mux_right_track_16.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _951_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_279_),
    .Z(\mux_right_track_16.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _952_ (.A(\mux_bottom_track_17.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_280_),
    .Z(\mux_bottom_track_17.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _953_ (.A(\mux_bottom_track_17.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_281_),
    .Z(\mux_bottom_track_17.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _954_ (.A(\mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_282_),
    .Z(\mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _955_ (.A(net93),
    .TE_B(_283_),
    .Z(\mux_bottom_track_17.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _955__93 (.HI(net93));
 sky130_fd_sc_hd__ebufn_1 _956_ (.A(\mux_bottom_track_17.INVTX1_6_.out ),
    .TE_B(_284_),
    .Z(\mux_bottom_track_17.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _957_ (.A(\mux_bottom_track_17.INVTX1_4_.out ),
    .TE_B(_285_),
    .Z(\mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _958_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_286_),
    .Z(\mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _959_ (.A(\mux_bottom_track_17.INVTX1_1_.out ),
    .TE_B(_287_),
    .Z(\mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _960_ (.A(\mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_288_),
    .Z(\mux_bottom_track_17.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _961_ (.A(\mux_bottom_track_17.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_289_),
    .Z(\mux_bottom_track_17.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _962_ (.A(\mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_290_),
    .Z(\mux_bottom_track_17.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _963_ (.A(\mux_bottom_track_17.INVTX1_7_.out ),
    .TE_B(_291_),
    .Z(\mux_bottom_track_17.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _964_ (.A(\mux_bottom_track_17.INVTX1_5_.out ),
    .TE_B(_292_),
    .Z(\mux_bottom_track_17.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _965_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_293_),
    .Z(\mux_bottom_track_17.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _966_ (.A(\mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_294_),
    .Z(\mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _967_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_295_),
    .Z(\mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _968_ (.A(\mux_left_track_17.mux_l3_in_1_.TGATE_0_.out ),
    .TE_B(_296_),
    .Z(\mux_left_track_17.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _969_ (.A(\mux_left_track_17.mux_l2_in_3_.TGATE_0_.out ),
    .TE_B(_297_),
    .Z(\mux_left_track_17.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _970_ (.A(\mux_left_track_17.mux_l2_in_1_.TGATE_0_.out ),
    .TE_B(_298_),
    .Z(\mux_left_track_17.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _971_ (.A(net94),
    .TE_B(_299_),
    .Z(\mux_left_track_17.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__conb_1 _971__94 (.HI(net94));
 sky130_fd_sc_hd__ebufn_1 _972_ (.A(\mux_left_track_17.INVTX1_6_.out ),
    .TE_B(_300_),
    .Z(\mux_left_track_17.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _973_ (.A(\mux_bottom_track_17.INVTX1_3_.out ),
    .TE_B(_301_),
    .Z(\mux_left_track_17.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _974_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_302_),
    .Z(\mux_left_track_17.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _975_ (.A(\mux_bottom_track_9.INVTX1_1_.out ),
    .TE_B(_303_),
    .Z(\mux_left_track_17.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_2 _976_ (.A(\mux_left_track_17.mux_l3_in_0_.TGATE_0_.out ),
    .TE_B(_304_),
    .Z(\mux_left_track_17.mux_l4_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _977_ (.A(\mux_left_track_17.mux_l2_in_2_.TGATE_0_.out ),
    .TE_B(_305_),
    .Z(\mux_left_track_17.mux_l3_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _978_ (.A(\mux_left_track_17.mux_l2_in_0_.TGATE_0_.out ),
    .TE_B(_306_),
    .Z(\mux_left_track_17.mux_l3_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _979_ (.A(\mux_left_track_17.INVTX1_7_.out ),
    .TE_B(_307_),
    .Z(\mux_left_track_17.mux_l2_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _980_ (.A(\mux_left_track_17.INVTX1_5_.out ),
    .TE_B(_308_),
    .Z(\mux_left_track_17.mux_l2_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _981_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_309_),
    .Z(\mux_left_track_17.mux_l2_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _982_ (.A(\mux_left_track_17.mux_l1_in_0_.TGATE_0_.out ),
    .TE_B(_310_),
    .Z(\mux_left_track_17.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 _983_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_311_),
    .Z(\mux_left_track_17.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_2_0__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_2_1__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_2_2__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_2_3__leaf_prog_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\mem_bottom_track_1.DFF_0_.D ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\mem_top_track_16.DFF_0_.D ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\mem_bottom_track_17.DFF_3_.Q ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\mem_top_track_0.DFF_3_.Q ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\mem_left_track_17.DFF_0_.Q ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\mem_left_track_1.DFF_3_.Q ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\mem_left_track_1.DFF_0_.Q ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\mem_top_track_8.DFF_0_.Q ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\mem_bottom_track_1.DFF_0_.Q ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\mem_bottom_track_17.DFF_0_.Q ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\mem_right_track_8.DFF_0_.Q ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\mem_right_track_0.DFF_0_.D ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\mem_right_track_16.DFF_2_.Q ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\mem_bottom_track_9.DFF_2_.Q ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\mem_right_track_8.DFF_2_.Q ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\mem_right_track_0.DFF_2_.Q ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\mem_top_track_0.DFF_2_.Q ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\mem_bottom_track_1.DFF_2_.Q ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\mem_left_track_9.DFF_0_.Q ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\mem_left_track_1.DFF_2_.Q ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\mem_left_track_9.DFF_2_.Q ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\mem_bottom_track_9.DFF_1_.Q ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\mem_top_track_16.DFF_0_.Q ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\mem_left_track_17.DFF_2_.Q ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\mem_top_track_16.DFF_2_.Q ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\mem_top_track_0.DFF_0_.Q ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\mem_top_track_8.DFF_2_.Q ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\mem_right_track_0.DFF_0_.Q ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\mem_bottom_track_17.DFF_2_.Q ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\mem_bottom_track_9.DFF_0_.Q ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\mem_right_track_0.DFF_1_.Q ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\mem_right_track_8.DFF_1_.Q ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mem_left_track_1.DFF_1_.Q ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\mem_bottom_track_1.DFF_3_.Q ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\mem_bottom_track_17.DFF_1_.Q ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\mem_top_track_8.DFF_1_.Q ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\mem_left_track_17.DFF_1_.Q ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\mem_bottom_track_1.DFF_1_.Q ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\mem_top_track_16.DFF_1_.Q ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\mem_top_track_0.DFF_1_.Q ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\mem_left_track_9.DFF_1_.Q ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mem_right_track_16.DFF_1_.Q ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\mem_left_track_17.DFF_0_.D ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\mem_right_track_16.DFF_0_.Q ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\mem_right_track_16.DFF_0_.D ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\mem_bottom_track_17.DFF_0_.D ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\mem_right_track_0.DFF_3_.Q ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(chanx_left_in[6]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(chanx_left_in[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(chanx_left_in[8]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(chanx_right_in[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(chanx_right_in[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(chanx_right_in[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(chanx_right_in[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chanx_right_in[4]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(chanx_right_in[5]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(chanx_right_in[6]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(chanx_right_in[7]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(chanx_right_in[8]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(chany_bottom_in[0]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(chany_bottom_in[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chany_bottom_in[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chany_bottom_in[3]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(chany_bottom_in[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(chany_bottom_in[5]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(chany_bottom_in[6]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(chany_bottom_in[7]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ccff_head),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(chany_bottom_in[8]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(chany_top_in[0]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(chany_top_in[1]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(chany_top_in[2]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(chany_top_in[3]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(chany_top_in[4]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(chany_top_in[5]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(chany_top_in[6]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(chany_top_in[7]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(chany_top_in[8]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(chanx_left_in[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(chanx_left_in[1]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(chanx_left_in[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(chanx_left_in[3]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(chanx_left_in[4]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(chanx_left_in[5]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(ccff_tail));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output53 (.A(net53),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(chany_top_out[8]));
endmodule

